library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_signed.all ;
use ieee.std_logic_arith.all;
library work;
use work.pkg2.all;

package pkg2 is
  type Arr_type is array (0 to 12) of std_logic_vector(13 downto 0);
end package;

package body pkg2 is
end package body;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_signed.all ;
use ieee.std_logic_arith.all;
library work;
use work.pkg2.all;

entity noteTable is
port(
  CLK     					: in std_logic;
  resetN 					: in std_logic;
  addrArr    				: in Arr_type;
  sound_choose				: in std_logic_vector(1 downto 0);
  Q       					: out std_logic_vector(15 downto 0)
);
end noteTable;

architecture arch of noteTable is
	constant array_size 			: integer := 8201 ;

	type table_type is array(0 to array_size - 1) of std_logic_vector(15 downto 0);
	signal arr_table				: table_type;
	signal Q_tmp       			:  std_logic_vector(15 downto 0) ;
	constant sound0 : table_type := (X"0008",X"FFF8",X"0006",X"FFFF",X"0000",X"0007",X"FFFF",X"FFF7",X"0007",X"0006",X"FFF4",X"FFF4",X"FFF8",X"FFFB",X"0000",X"FFF8",X"FFF7",X"FFF9",X"FFFE",X"FFFF",X"FFFF",X"0000",X"0004",X"FFFB",X"0008",X"FFFF",X"0004",X"FFFC",X"FFFD",X"0000",X"0008",X"0004",X"000A",X"0007",X"000F",X"0001",X"FFF5",X"0002",X"0002",X"FFFB",X"0000",X"0000",X"0005",X"0001",X"FFF4",X"0000",X"FFF4",X"FFF2",X"FFFD",X"FFF9",X"FFF7",X"0004",X"0005",X"0002",X"0004",X"FFFE",X"0006",X"0000",X"0007",X"0009",X"0001",X"0002",X"0005",X"0008",X"FFFE",X"FFF8",X"FFF7",X"0000",X"FFF7",X"FFFA",X"0004",X"0003",X"0001",X"FFFE",X"0006",X"FFFC",X"0002",X"000D",X"FFFC",X"0002",X"FFF9",X"0000",X"0000",X"FFFF",X"0005",X"0001",X"FFFF",X"FFF8",X"0000",X"FFFF",X"FFEE",X"FFF6",X"FFF2",X"0002",X"FFFF",X"FFFD",X"FFFB",X"0001",X"0008",X"0006",X"0005",X"0004",X"0000",X"FFF5",X"0007",X"0009",X"FFFB",X"0000",X"0008",X"0000",X"FFF9",X"0000",X"FFF7",X"0000",X"0000",X"FFFE",X"0000",X"FFF7",X"FFF8",X"FFFC",X"0001",X"FFFE",X"FFF6",X"FFFB",X"FFFB",X"FFFA",X"FFF8",X"FFF0",X"FFFC",X"0000",X"000B",X"000F",X"0004",X"0000",X"0001",X"FFFC",X"000E",X"FFF7",X"FFF9",X"0005",X"FFFB",X"0003",X"0001",X"FFF8",X"FFF8",X"FFF7",X"FFF9",X"FFF9",X"FFFA",X"0001",X"0000",X"0003",X"0000",X"FFFF",X"0000",X"0004",X"FFF8",X"0008",X"0005",X"FFF8",X"0004",X"FFFC",X"0004",X"FFFA",X"FFFA",X"0001",X"FFFE",X"0007",X"0000",X"0003",X"0000",X"0001",X"FFFE",X"FFF7",X"FFF0",X"0000",X"0007",X"0002",X"FFFB",X"0000",X"0008",X"0002",X"FFFC",X"FFFE",X"FFFD",X"0002",X"0003",X"0002",X"FFFB",X"0003",X"0001",X"0003",X"0000",X"000B",X"FFF8",X"FFF5",X"0004",X"000B",X"0006",X"0003",X"FFFB",X"FFF1",X"FFFF",X"0010",X"FFFE",X"0005",X"FFF8",X"FFF6",X"FFFE",X"0000",X"0008",X"FFFB",X"0004",X"0000",X"0001",X"FFFF",X"FFFA",X"0000",X"FFF5",X"FFFB",X"0001",X"FFF8",X"FFFD",X"FFFC",X"000F",X"FFFF",X"FFFF",X"0000",X"FFFD",X"0002",X"0000",X"0004",X"0000",X"FFFA",X"FFFD",X"FFFA",X"000B",X"0008",X"0007",X"000E",X"0000",X"FFF6",X"0000",X"0007",X"FFFE",X"0004",X"FFFB",X"FFFE",X"FFF7",X"FFF9",X"FFFE",X"0006",X"0007",X"FFFF",X"0000",X"FFF6",X"0000",X"FFFD",X"0003",X"0001",X"0008",X"0003",X"FFF9",X"000A",X"0009",X"000B",X"0007",X"0008",X"0003",X"FFF8",X"FFF8",X"FFF5",X"FFFE",X"0008",X"FFF6",X"0001",X"0001",X"FFF9",X"FFFB",X"FFFD",X"0000",X"0003",X"0000",X"0000",X"0002",X"0001",X"FFFF",X"0009",X"0005",X"FFFC",X"FFF9",X"FFF3",X"0001",X"FFFF",X"FFF6",X"FFED",X"FFF5",X"FFFD",X"0003",X"000E",X"FFFA",X"0007",X"FFFA",X"0000",X"0009",X"0000",X"0000",X"FFF3",X"FFFA",X"FFF1",X"0002",X"FFF6",X"FFFD",X"FFFE",X"FFFA",X"0002",X"0003",X"0005",X"FFFD",X"FFFE",X"FFFF",X"0000",X"0001",X"FFFB",X"FFFD",X"0001",X"0001",X"0004",X"FFF8",X"0000",X"0014",X"000B",X"000C",X"FFF9",X"FFFE",X"0004",X"FFFF",X"0000",X"0006",X"0005",X"0000",X"FFFA",X"FFFB",X"000C",X"0001",X"FFFD",X"0000",X"0006",X"000A",X"FFFF",X"FFFD",X"0004",X"0001",X"0008",X"0000",X"FFFB",X"FFF3",X"FFFF",X"FFF4",X"FFEF",X"0006",X"0000",X"0005",X"0006",X"FFFF",X"FFFE",X"0001",X"000B",X"0005",X"FFFF",X"0000",X"FFFE",X"FFF7",X"FFF8",X"FFFD",X"0003",X"0005",X"0005",X"0000",X"FFF7",X"FFF6",X"FFF4",X"0006",X"0000",X"0002",X"0003",X"FFFE",X"FFFD",X"FFF6",X"0001",X"0006",X"0004",X"FFFE",X"0000",X"FFFE",X"0004",X"0007",X"0001",X"FFFC",X"FFFF",X"0002",X"0004",X"FFF9",X"0005",X"0005",X"0000",X"0001",X"FFFD",X"FFFE",X"0000",X"0001",X"FFF6",X"FFFC",X"0007",X"FFFE",X"0000",X"000A",X"0002",X"0002",X"0000",X"0001",X"FFF8",X"FFFD",X"0007",X"FFF2",X"FFF7",X"FFF7",X"FFFB",X"FFFA",X"0001",X"0000",X"0002",X"0009",X"FFFC",X"0004",X"0007",X"0004",X"0009",X"FFFA",X"0003",X"FFF8",X"0001",X"0003",X"0004",X"0008",X"0000",X"000C",X"0004",X"FFFE",X"FFF9",X"FFFB",X"0000",X"0001",X"FFFC",X"0001",X"FFF9",X"FFF7",X"0004",X"0001",X"0000",X"0009",X"FFFD",X"FFF5",X"FFF9",X"FFF8",X"0002",X"0000",X"FFFE",X"000C",X"000A",X"0003",X"FFFE",X"FFFC",X"0000",X"0004",X"0003",X"0000",X"0002",X"FFFE",X"FFF2",X"FFFF",X"000B",X"0007",X"FFFE",X"FFFE",X"FFFF",X"0007",X"0004",X"0007",X"0001",X"FFF3",X"FFEF",X"FFFC",X"FFFB",X"FFFE",X"FFF5",X"0004",X"FFF3",X"0001",X"0007",X"0002",X"0008",X"000C",X"000C",X"0008",X"0009",X"000C",X"0002",X"FFF8",X"0000",X"0001",X"FFF8",X"FFF9",X"FFF1",X"FFF8",X"FFF8",X"FFFD",X"FFFC",X"0003",X"FFFD",X"FFF9",X"0005",X"0000",X"FFF4",X"FFF5",X"0003",X"000F",X"0007",X"000C",X"0005",X"0001",X"0006",X"FFFB",X"FFF9",X"0000",X"FFFB",X"0000",X"0003",X"000A",X"0000",X"FFF9",X"0001",X"0002",X"FFFC",X"FFFD",X"0001",X"0009",X"FFF4",X"FFEF",X"FFF7",X"0009",X"0006",X"0017",X"0001",X"FFFE",X"0007",X"FFFE",X"000C",X"0005",X"0003",X"0003",X"FFFA",X"FFF5",X"FFF1",X"000B",X"0001",X"FFF5",X"000D",X"0001",X"0008",X"FFFD",X"0006",X"FFF8",X"FFF0",X"FFED",X"FFFB",X"FFF2",X"0000",X"0002",X"0005",X"0009",X"0003",X"FFFC",X"0006",X"0007",X"FFFD",X"0009",X"000B",X"0007",X"FFF2",X"FFFE",X"FFF7",X"FFFB",X"FFFE",X"FFF9",X"FFFA",X"0009",X"FFFE",X"FFF4",X"0005",X"0007",X"0000",X"FFFE",X"000B",X"0009",X"FFF9",X"FFF4",X"0003",X"FFF3",X"FFEA",X"FFF4",X"FFFE",X"0007",X"0007",X"0012",X"000E",X"0003",X"FFF8",X"0010",X"000A",X"FFF8",X"FFFB",X"0008",X"FFF9",X"FFED",X"FFF9",X"FFF2",X"0009",X"FFFB",X"000C",X"0019",X"0004",X"0002",X"0000",X"FFF8",X"0000",X"0009",X"FFF9",X"0005",X"0010",X"0000",X"0003",X"0004",X"0006",X"FFEE",X"FFFD",X"0004",X"FFF6",X"FFF1",X"0002",X"0005",X"0000",X"FFF3",X"0004",X"0015",X"0005",X"0002",X"000B",X"0007",X"0000",X"FFFC",X"0004",X"0003",X"FFF0",X"FFFB",X"0004",X"FFF5",X"FFFB",X"FFFC",X"0005",X"0000",X"000E",X"0018",X"000C",X"000C",X"FFF6",X"FFFA",X"FFFD",X"FFF6",X"FFFE",X"0008",X"0002",X"FFFF",X"FFFD",X"FFFE",X"0003",X"FFFE",X"0004",X"0011",X"0011",X"0003",X"FFFD",X"FFFC",X"FFF8",X"FFF6",X"0001",X"000B",X"FFE8",X"FFF2",X"FFFD",X"FFE1",X"FFDB",X"FFEB",X"FFF4",X"FFE6",X"FFEE",X"0006",X"0002",X"FFFD",X"002B",X"0029",X"002C",X"003F",X"0041",X"004A",X"003A",X"0057",X"004A",X"004F",X"0036",X"FEFD",X"FEA2",X"FFB9",X"FFFC",X"0024",X"FF92",X"FEC2",X"0166",X"0395",X"0310",X"0312",X"010D",X"00E1",X"FE2D",X"FA0C",X"F3E5",X"F06A",X"F607",X"F896",X"00B6",X"0E2F",X"1832",X"1B6E",X"1848",X"0F7A",X"FB61",X"EC13",X"E59D",X"E7EE",X"F1A2",X"F7CC",X"FCB5",X"0231",X"0B70",X"0DD0",X"0A94",X"0CDD",X"0BC6",X"0370",X"023C",X"02E3",X"FAF3",X"F0C3",X"E59D",X"E361",X"EFA3",X"F7FE",X"FFA3",X"09DA",X"18B1",X"1FED",X"1A52",X"1AD4",X"1A28",X"0889",X"F2F5",X"EE3C",X"ECE0",X"EA51",X"E211",X"D6C0",X"E186",X"F48A",X"067B",X"16E1",X"253B",X"2B34",X"2025",X"0FBA",X"052A",X"FE05",X"F178",X"EB63",X"F14F",X"F8A7",X"FA73",X"EAB5",X"E00E",X"E5A6",X"F215",X"01D5",X"174D",X"2B1C",X"2FDB",X"27EA",X"1C1B",X"0D82",X"F6CE",X"E1DA",X"E040",X"E661",X"EDDE",X"E68F",X"DA87",X"E6E7",X"FD87",X"0C5C",X"19E6",X"2C54",X"35C1",X"2A3D",X"146A",X"FE54",X"ED1F",X"DBE2",X"D82E",X"E704",X"FC88",X"031C",X"F06F",X"E918",X"F853",X"0476",X"073D",X"0F47",X"1E0A",X"22C0",X"1C30",X"0E90",X"008D",X"F491",X"EE53",X"F3B1",X"FCA1",X"0077",X"EEEE",X"DCB6",X"E7D9",X"FD25",X"02F9",X"040F",X"0F03",X"18DE",X"19CA",X"14BF",X"0C75",X"03F3",X"F841",X"F4D0",X"F8C0",X"FF3B",X"F661",X"DDC5",X"D878",X"EEB3",X"0287",X"066A",X"0D8C",X"1AC6",X"1F84",X"1BAE",X"1302",X"0B20",X"FF5F",X"F6FC",X"F3CE",X"F6A1",X"F98D",X"E85B",X"D5C5",X"E21A",X"FE13",X"09DB",X"0AEA",X"1346",X"17F0",X"170C",X"11FC",X"0A48",X"FF95",X"F7AC",X"F85B",X"FD41",X"072F",X"01E0",X"E7AD",X"DD04",X"EE38",X"FCB5",X"FB03",X"FFFE",X"0BA3",X"12D3",X"1597",X"13B0",X"0C4C",X"0067",X"FB30",X"FAB9",X"033E",X"0C04",X"FD18",X"E400",X"E3B1",X"F54A",X"F9AE",X"F875",X"0100",X"09AB",X"1068",X"139D",X"1434",X"0CFD",X"04B2",X"FDD0",X"FC2B",X"0835",X"0881",X"EDDF",X"D937",X"E1A5",X"EE10",X"F048",X"FBEA",X"0BDF",X"1832",X"1D0D",X"1E1B",X"1963",X"0D71",X"0003",X"F1C5",X"F43E",X"0315",X"FC17",X"E5B2",X"E42A",X"F584",X"F956",X"F86C",X"FEEA",X"07AD",X"0E8A",X"11B4",X"135B",X"0DBB",X"0719",X"FDF0",X"F9A6",X"0922",X"1153",X"FBF4",X"E4DE",X"E79D",X"ED9A",X"EB35",X"F0C4",X"FD39",X"0B13",X"126F",X"17AB",X"1578",X"0EC6",X"066E",X"F9E5",X"FDE0",X"1058",X"0C88",X"F138",X"E4A0",X"EBDB",X"EC8F",X"ECEF",X"F3F1",X"01A7",X"0D75",X"15D0",X"192E",X"14B9",X"0ED3",X"0277",X"F995",X"069D",X"1196",X"FE2C",X"E245",X"DFD3",X"E4C0",X"E574",X"EADF",X"F912",X"0AF7",X"187F",X"224A",X"219D",X"1AFE",X"0F2E",X"FC92",X"FA23",X"0A06",X"09A8",X"EED9",X"DEDB",X"E2E3",X"E5D8",X"E7FE",X"EF28",X"FEDE",X"0C70",X"1803",X"1D6B",X"19DF",X"1459",X"0631",X"F99A",X"0390",X"1213",X"0536",X"EB7F",X"E5F1",X"E89E",X"EA53",X"EC9E",X"F5F3",X"01A6",X"0C62",X"1675",X"1730",X"1477",X"0D47",X"FD31",X"FAB4",X"0D08",X"1287",X"F9CE",X"E6A4",X"E3F6",X"E5B7",X"E7CE",X"EF73",X"FDA6",X"0A3E",X"1700",X"1D2E",X"1C05",X"19B1",X"0BCE",X"FB22",X"FFBB",X"0F1A",X"0439",X"EA35",X"DECB",X"DD80",X"DEF9",X"E389",X"F110",X"01C0",X"1325",X"2282",X"2578",X"239C",X"1AE3",X"05D6",X"F984",X"04D0",X"098A",X"F2FD",X"DF37",X"DAC9",X"DF08",X"E51A",X"F137",X"01BC",X"108E",X"1ED5",X"2323",X"1EC8",X"193E",X"089C",X"F2DF",X"F281",X"0461",X"00C9",X"EE01",X"E40C",X"E665",X"EBE4",X"F227",X"FCEF",X"078A",X"130F",X"1C03",X"1ACC",X"17C5",X"1010",X"FBAC",X"ECC4",X"FAA7",X"082F",X"FD98",X"ED62",X"E7A3",X"EA9E",X"EE52",X"F510",X"FE4B",X"08DE",X"15F2",X"1B29",X"193D",X"16EE",X"0A42",X"F32A",X"F0C3",X"0468",X"0803",X"F9A1",X"ED81",X"EC1A",X"ED86",X"EF6A",X"F500",X"FB8F",X"06CC",X"1226",X"14F2",X"16E9",X"156A",X"048F",X"F370",X"FE89",X"0D27",X"072F",X"F70A",X"EE39",X"EC89",X"EADC",X"ED50",X"F29A",X"FB9F",X"0A8A",X"13D3",X"1739",X"1A8E",X"1468",X"FD8C",X"F6B5",X"054C",X"0A1E",X"FCBC",X"EE3F",X"EA74",X"EA32",X"EC48",X"F207",X"F8CC",X"0554",X"11E7",X"1692",X"18A4",X"1A7B",X"0A59",X"F5E2",X"FB38",X"085C",X"049F",X"F426",X"EA1F",X"E8BD",X"E9CD",X"EF96",X"F5DC",X"FE50",X"0BFA",X"1537",X"17E2",X"1C5E",X"1810",X"00E2",X"F5C2",X"00E7",X"0826",X"FD95",X"EEA9",X"E98F",X"E97F",X"EC60",X"F158",X"F5D5",X"00E4",X"0DC1",X"142E",X"18CB",X"1EDC",X"1107",X"FAA7",X"FA6F",X"0770",X"0802",X"F92F",X"ED4B",X"E940",X"E827",X"EBA8",X"EF3D",X"F7B8",X"068B",X"12B1",X"1739",X"1F3D",X"1E8E",X"0772",X"F719",X"FDDA",X"07CD",X"0092",X"F166",X"E977",X"E71C",X"EA3C",X"EF46",X"F470",X"FFB4",X"0E4A",X"14CC",X"1933",X"2143",X"158E",X"FDB6",X"F74C",X"0297",X"066B",X"F9D4",X"ED84",X"E8B4",X"E912",X"ED34",X"EFC7",X"F5EC",X"03A6",X"100B",X"14BA",X"1EB7",X"212B",X"0D7B",X"FA68",X"FC93",X"06C8",X"036C",X"F5FC",X"ECE0",X"E899",X"E9EB",X"EBD4",X"EE90",X"F810",X"07EE",X"100D",X"1727",X"2202",X"1AA7",X"03AF",X"F8A8",X"019E",X"0863",X"FF58",X"F375",X"EC01",X"EB2C",X"EDC5",X"EFB5",X"F2BF",X"FE78",X"0A22",X"0E79",X"1973",X"1FC9",X"10F2",X"FCA2",X"FAFB",X"062E",X"066B",X"FB70",X"F106",X"EBF9",X"EC76",X"EE6A",X"EF1B",X"F523",X"0313",X"0A25",X"11D3",X"1F51",X"1E3B",X"09E6",X"FADC",X"FF84",X"06E6",X"0116",X"F5B2",X"ED07",X"EB25",X"ED0A",X"EEBF",X"F06B",X"FC22",X"07DB",X"0CC4",X"17EF",X"214D",X"15FA",X"FFE3",X"F8D4",X"02BA",X"063F",X"FEEE",X"F469",X"EE4E",X"ED6C",X"EF77",X"EF0C",X"F3BB",X"00B7",X"0761",X"0DBE",X"1B3E",X"1DFD",X"0C24",X"FA3D",X"FCE6",X"05A8",X"046A",X"FB0C",X"F220",X"EE76",X"F031",X"F16A",X"F0D3",X"FA51",X"0428",X"0719",X"1051",X"1CA2",X"1721",X"01CB",X"F8AF",X"008D",X"0699",X"02A4",X"F932",X"F227",X"F0AE",X"F2E3",X"F019",X"F1F8",X"FCC3",X"02A9",X"076C",X"159D",X"1D7E",X"0FB0",X"FD19",X"FCD7",X"05F5",X"0881",X"012A",X"F74E",X"F082",X"F07E",X"EF61",X"EC5D",X"F411",X"FEA5",X"02CB",X"0CDD",X"1C31",X"1C37",X"089B",X"FC6A",X"0119",X"0821",X"05DA",X"FC4C",X"F296",X"EF06",X"F079",X"ECC4",X"EDEE",X"F8EE",X"FFBC",X"04D3",X"135A",X"1F90",X"15A2",X"0286",X"FD9E",X"04CD",X"089C",X"02FE",X"F946",X"F11E",X"F15F",X"F04C",X"EC62",X"F251",X"FBDF",X"FFC5",X"0823",X"18A3",X"1CAE",X"0BE3",X"FD2D",X"FEFC",X"07B2",X"08CF",X"0211",X"F76E",X"F232",X"F1E0",X"ED01",X"EC77",X"F5C4",X"FC22",X"003E",X"0DAC",X"1D01",X"181F",X"05F9",X"FD9E",X"0398",X"0915",X"0673",X"FD33",X"F3E8",X"F28C",X"F068",X"EAF5",X"EF6F",X"F90E",X"FCBB",X"033A",X"1546",X"1ED0",X"1278",X"01EE",X"FFF3",X"073C",X"098C",X"0420",X"F864",X"F23E",X"F1DB",X"EC1B",X"E9C7",X"F250",X"F9D2",X"FC88",X"093B",X"1BC5",X"1C9D",X"0C19",X"0041",X"0322",X"0868",X"089B",X"FFFB",X"F5AE",X"F36F",X"F0D3",X"EA4F",X"ECE9",X"F6A1",X"FA68",X"FF09",X"10A1",X"1E27",X"1691",X"0584",X"0062",X"04CE",X"08C7",X"05AE",X"FAA9",X"F439",X"F3B4",X"EE3E",X"EA70",X"F159",X"F8B1",X"FA49",X"04FD",X"184E",X"1E5F",X"10E9",X"034D",X"0231",X"067E",X"0824",X"0050",X"F574",X"F31C",X"F0DA",X"EA6C",X"EBAE",X"F593",X"FA0F",X"FDD5",X"0E22",X"1E4A",X"1B31",X"0A67",X"0197",X"02EC",X"076C",X"0632",X"FBD4",X"F516",X"F3FC",X"EE82",X"E93F",X"EF06",X"F730",X"F906",X"01DC",X"14EA",X"1F34",X"1469",X"05E3",X"01A8",X"050C",X"08E1",X"0354",X"F947",X"F5F6",X"F34B",X"EBD3",X"EAFA",X"F3E0",X"F7E3",X"F9C4",X"070B",X"19A3",X"1B5F",X"0D8B",X"0307",X"01EF",X"06DC",X"07AE",X"FEA7",X"F74F",X"F597",X"F080",X"EA91",X"EF46",X"F720",X"F880",X"FE82",X"10C3",X"1E8D",X"1811",X"0978",X"011F",X"01F8",X"0657",X"023B",X"F902",X"F5A1",X"F461",X"EDF4",X"EBF7",X"F3E1",X"F88A",X"F9AA",X"0471",X"17C5",X"1D12",X"112A",X"041F",X"FF6A",X"041E",X"073E",X"00F2",X"FA50",X"F8EE",X"F43B",X"EC37",X"EE12",X"F4C5",X"F632",X"F8CC",X"0910",X"1991",X"17F1",X"0B72",X"019D",X"01DC",X"0827",X"0731",X"FF67",X"FB8C",X"F9E2",X"F1C1",X"ECAD",X"F13E",X"F573",X"F432",X"FBB6",X"0F09",X"1955",X"1354",X"0790",X"0118",X"04D9",X"090C",X"03F7",X"FCF1",X"FB4A",X"F6BA",X"EE11",X"ED9E",X"F3B4",X"F4FF",X"F543",X"0387",X"15F9",X"19BC",X"106D",X"049C",X"01D6",X"06E0",X"06DB",X"0009",X"FBEF",X"FA7B",X"F26C",X"EC0A",X"EF31",X"F440",X"F2D9",X"F85B",X"0B50",X"18F9",X"175B",X"0BE7",X"0318",X"0509",X"096B",X"05B7",X"FEA3",X"FD0C",X"F86A",X"EF3F",X"EC4D",X"F191",X"F317",X"F1B8",X"FDA6",X"10B4",X"18F7",X"12E4",X"0701",X"02AD",X"074B",X"0907",X"02CA",X"FEB1",X"FCDF",X"F588",X"EDAD",X"EED4",X"F3DD",X"F216",X"F4BB",X"0510",X"14B6",X"1750",X"0E10",X"0426",X"045F",X"092D",X"06C5",X"006C",X"FE7B",X"FA91",X"F17C",X"EC9B",X"F0CC",X"F2A1",X"F025",X"F947",X"0BC0",X"17C4",X"15EA",X"0B10",X"04CF",X"07D6",X"09E8",X"03EF",X"FF83",X"FD7E",X"F6C0",X"ED90",X"ECF1",X"F1F3",X"F02A",X"F176",X"FFFE",X"11A9",X"18FB",X"1273",X"07E0",X"0549",X"09A0",X"07A8",X"01CA",X"FF7C",X"FC6F",X"F396",X"ECE5",X"F06F",X"F23F",X"EF29",X"F554",X"066D",X"1518",X"16DC",X"0D4D",X"04BF",X"06B7",X"096B",X"04B1",X"0042",X"FEB4",X"F979",X"EFD6",X"EE4B",X"F32E",X"F1CE",X"F0F5",X"FC1B",X"0D78",X"1805",X"1494",X"0968",X"0489",X"07E1",X"0688",X"00EA",X"FE62",X"FCEF",X"F584",X"EE73",X"F18E",X"F40A",X"F0D1",X"F41B",X"0270",X"1294",X"17BA",X"0FCD",X"057D",X"054C",X"07E5",X"048C",X"00C5",X"0025",X"FCC3",X"F2F4",X"EFAC",X"F32F",X"F186",X"EF02",X"F696",X"077A",X"14BE",X"152E",X"0AE8",X"04FE",X"07C3",X"07AF",X"0365",X"00F6",X"0088",X"F968",X"F147",X"F282",X"F453",X"F0A5",X"F0B9",X"FC38",X"0C9A",X"1583",X"1059",X"0626",X"04E0",X"079A",X"059B",X"01B1",X"01A2",X"FF2B",X"F5BE",X"F163",X"F44F",X"F38F",X"F012",X"F440",X"02EA",X"11B6",X"1585",X"0C6C",X"0526",X"0644",X"06E7",X"035A",X"0130",X"01AE",X"FB98",X"F2F2",X"F293",X"F454",X"F142",X"EF59",X"F7F7",X"07EE",X"142C",X"1275",X"08F2",X"05E8",X"07AA",X"06C6",X"0313",X"0360",X"01E9",X"F8DF",X"F2EE",X"F3F3",X"F335",X"EE80",X"EFE5",X"FC12",X"0C69",X"13FC",X"0D90",X"0683",X"0686",X"087D",X"05AA",X"03CC",X"04E3",X"FF7D",X"F649",X"F388",X"F47B",X"F0FF",X"ED5C",X"F2C6",X"01D7",X"10E5",X"129D",X"0AC7",X"067A",X"0824",X"07B8",X"03E8",X"0427",X"034A",X"FAE1",X"F3DA",X"F3CB",X"F396",X"EF40",X"EEDF",X"F887",X"0966",X"1416",X"104E",X"088E",X"0689",X"07ED",X"0517",X"030F",X"049A",X"006E",X"F7C7",X"F401",X"F4CE",X"F21A",X"EE16",X"F0AE",X"FDAE",X"0DF3",X"128C",X"0C6B",X"06EA",X"07D1",X"07E3",X"04B8",X"0581",X"0578",X"FE59",X"F669",X"F4E1",X"F418",X"EF73",X"ECF1",X"F305",X"036E",X"1048",X"104D",X"095C",X"06DA",X"08B6",X"069A",X"04FB",X"06AE",X"03B6",X"FAF4",X"F58C",X"F51B",X"F23F",X"EDB0",X"ED49",X"F84B",X"0969",X"1211",X"0E76",X"0899",X"08BE",X"08A0",X"0536",X"0566",X"0605",X"0005",X"F7C2",X"F514",X"F44A",X"F08B",X"ECB5",X"F031",X"FF5A",X"0E60",X"11D4",X"0BA6",X"07B7",X"0894",X"062E",X"0442",X"060B",X"04C9",X"FCFD",X"F6E0",X"F5F4",X"F3AE",X"EF14",X"EC58",X"F4E7",X"0592",X"10E8",X"0FA2",X"0950",X"0856",X"07E6",X"04D0",X"04B3",X"0636",X"01CD",X"F9B8",X"F698",X"F595",X"F2B6",X"ED9B",X"EE98",X"FB77",X"0BA4",X"1241",X"0D1F",X"0857",X"081E",X"05B5",X"033D",X"04C7",X"04A5",X"FDBE",X"F80A",X"F692",X"F592",X"F185",X"ED2C",X"F2B3",X"020E",X"0FC9",X"1115",X"0AC5",X"087E",X"075C",X"040A",X"0363",X"0578",X"029C",X"FB50",X"F78C",X"F679",X"F48B",X"EECE",X"ED38",X"F735",X"07B0",X"1183",X"0E97",X"09F7",X"08FA",X"066D",X"036D",X"0479",X"055E",X"FF87",X"F9CA",X"F734",X"F68E",X"F2A5",X"ED13",X"EFAC",X"FCF4",X"0C95",X"10DE",X"0C35",X"0966",X"07B5",X"03FF",X"0262",X"0524",X"0379",X"FDCC",X"F9B0",X"F8AC",X"F753",X"F159",X"ED56",X"F384",X"02D1",X"0EA6",X"0E38",X"09FC",X"0847",X"05B3",X"0257",X"03C3",X"059E",X"0213",X"FCA9",X"F97A",X"F8FB",X"F539",X"EEA8",X"EDD4",X"F854",X"0863",X"0F61",X"0CC0",X"09FA",X"081B",X"044B",X"0250",X"04DC",X"0452",X"FF8A",X"FA9A",X"F93F",X"F840",X"F2A1",X"ED4B",X"F078",X"FE97",X"0C20",X"0E8A",X"0BAB",X"09CC",X"0752",X"0346",X"03F1",X"0577",X"02F1",X"FD90",X"F9BA",X"F961",X"F65D",X"EFE8",X"EC91",X"F44D",X"0413",X"0D67",X"0D54",X"0B05",X"096A",X"0525",X"02D9",X"04D4",X"0560",X"01E3",X"FC7F",X"FA82",X"F972",X"F468",X"EDA7",X"ED93",X"F9A0",X"080C",X"0D31",X"0BF0",X"0AB2",X"07EA",X"0387",X"0394",X"05A9",X"04F8",X"0008",X"FBAB",X"FAC5",X"F838",X"F1BA",X"EC31",X"F0D2",X"FF7A",X"0A7E",X"0C91",X"0B4D",X"0A2A",X"05B4",X"02F2",X"046A",X"05FD",X"03AA",X"FE24",X"FB7E",X"FA59",X"F610",X"EEF9",X"EC2E",X"F5EF",X"0465",X"0BF0",X"0C1C",X"0BB5",X"08CA",X"0422",X"035C",X"0545",X"05D2",X"0173",X"FCD1",X"FB5D",X"F957",X"F3C7",X"EC9A",X"EE59",X"FB02",X"079B",X"0BE2",X"0C2D",X"0B5F",X"06DB",X"0392",X"0402",X"063C",X"04B7",X"FF85",X"FC69",X"FB21",X"F7E2",X"F0AA",X"EB9A",X"F210",X"FFE3",X"0941",X"0BA0",X"0C71",X"0A10",X"059C",X"03BB",X"0531",X"066D",X"02B8",X"FE20",X"FC2C",X"FA79",X"F5A1",X"ED88",X"EC80",X"F6D5",X"042A",X"0A60",X"0C63",X"0C5F",X"0874",X"04B8",X"03F7",X"0614",X"0522",X"0040",X"FD0B",X"FBB2",X"F9AC",X"F29B",X"EC28",X"EF92",X"FC75",X"06F8",X"0B03",X"0CD1",X"0AE5",X"06CD",X"03DD",X"04B3",X"0638",X"0322",X"FF05",X"FCCB",X"FBFD",X"F7EC",X"EFB5",X"EBDF",X"F39B",X"008F",X"0801",X"0BAB",X"0C64",X"099F",X"0571",X"03BC",X"05DD",X"05A9",X"01AA",X"FE37",X"FCF5",X"FBAF",X"F538",X"ED5A",X"ED67",X"F890",X"036D",X"0948",X"0C70",X"0BDC",X"0826",X"042D",X"044B",X"0634",X"03EF",X"0021",X"FD65",X"FD18",X"FA03",X"F23E",X"EC0E",X"F0DE",X"FCC1",X"0577",X"0ADA",X"0CBC",X"0AD8",X"0665",X"0395",X"0575",X"05A0",X"02A7",X"FEC4",X"FD75",X"FCAF",X"F7BE",X"EF4D",X"EC9A",X"F54B",X"FFBF",X"076E",X"0BFF",X"0C80",X"0968",X"04D6",X"0463",X"05DD",X"04BC",X"00E6",X"FDFE",X"FDB6",X"FBC5",X"F4F1",X"ED20",X"EF68",X"F947",X"0296",X"093D",X"0C4E",X"0BAC",X"0744",X"03E8",X"04E9",X"0555",X"0319",X"FF48",X"FE0B",X"FDD6",X"FA67",X"F1C8",X"ED38",X"F342",X"FCF8",X"0555",X"0ABD",X"0C81",X"0A28",X"0503",X"03E6",X"0502",X"04A9",X"013E",X"FE82",X"FE5B",X"FDB1",X"F7ED",X"EF41",X"EF14",X"F6C5",X"FFD6",X"0748",X"0B38",X"0BDC",X"0777",X"03E8",X"0425",X"0521",X"0399",X"002C",X"FEE0",X"FEF4",X"FD0A",X"F4AC",X"EE9C",X"F1B3",X"F9C3",X"0251",X"083A",X"0B99",X"0A2A",X"0595",X"03F7",X"0506",X"0579",X"0289",X"FFD8",X"FF00",X"FF46",X"FA55",X"F16A",X"EEB9",X"F3E9",X"FCA5",X"0499",X"09F8",X"0C25",X"0884",X"04B5",X"042A",X"0574",X"0433",X"010A",X"FEB0",X"FEE0",X"FE17",X"F6C0",X"EFBB",X"F074",X"F72C",X"0001",X"06CB",X"0BDB",X"0B2A",X"06C0",X"0403",X"04AB",X"0552",X"0304",X"0036",X"FED6",X"FFC5",X"FC13",X"F382",X"EF56",X"F242",X"FA65",X"0239",X"08D4",X"0C2A",X"0980",X"056B",X"0420",X"056A",X"0480",X"01EE",X"FF2B",X"FF68",X"FF51",X"F8B2",X"F13F",X"EF8F",X"F4C8",X"FCE6",X"044A",X"0A9F",X"0B9C",X"082A",X"04D4",X"0534",X"0572",X"03C9",X"00B9",X"FF0E",X"0045",X"FD9A",X"F5A0",X"F005",X"F0B5",X"F7C6",X"FF69",X"0716",X"0B9A",X"0A6E",X"065D",X"048E",X"0525",X"04B2",X"0293",X"FFC1",X"0018",X"00CC",X"FB32",X"F3A3",X"EF8C",X"F2FB",X"F9EE",X"0184",X"08AA",X"0B1E",X"0894",X"0538",X"0501",X"055D",X"0497",X"01D1",X"FFEE",X"016C",X"FF44",X"F839",X"F133",X"EFF3",X"F517",X"FC16",X"0447",X"0A36",X"0AF1",X"075F",X"0560",X"0579",X"0563",X"039C",X"0067",X"0081",X"0151",X"FCE6",X"F565",X"EFFA",X"F18F",X"F6FE",X"FE98",X"0686",X"0B28",X"09BF",X"0683",X"059C",X"05DA",X"0553",X"0242",X"FFE1",X"0136",X"FFEF",X"FA34",X"F2AB",X"EFFE",X"F31B",X"F967",X"01BB",X"0925",X"0B85",X"089C",X"0648",X"05C6",X"05DE",X"0465",X"0096",X"0069",X"0138",X"FE4F",X"F740",X"F0E7",X"F08D",X"F4A8",X"FC05",X"0498",X"0AD9",X"0A9B",X"07A5",X"0620",X"05E2",X"05ED",X"0299",X"000E",X"0110",X"00BD",X"FC44",X"F48A",X"F090",X"F1C7",X"F711",X"FED1",X"0754",X"0B1E",X"0932",X"06C5",X"05BC",X"061B",X"04BB",X"010C",X"00C0",X"01A2",X"0022",X"F992",X"F2E9",X"F0BD",X"F335",X"F92C",X"01D7",X"0927",X"0A77",X"0844",X"0666",X"05F5",X"064C",X"0304",X"00BA",X"0137",X"01A9",X"FE12",X"F6D0",X"F1C1",X"F12A",X"F4D8",X"FBFA",X"0501",X"0A33",X"099B",X"076F",X"05C9",X"067D",X"0547",X"01FB",X"011D",X"01D2",X"0128",X"FB81",X"F4AB",X"F0E3",X"F1CC",X"F67D",X"FEFB",X"0793",X"0A6D",X"0947",X"06DC",X"064A",X"06A9",X"0390",X"013F",X"0105",X"0214",X"FF6D",X"F925",X"F35B",X"F166",X"F351",X"F947",X"02AC",X"0921",X"09F8",X"07FA",X"05B7",X"0674",X"0503",X"0215",X"00A3",X"01CA",X"0202",X"FDC4",X"F723",X"F28B",X"F1CF",X"F4A9",X"FC60",X"0587",X"0991",X"0978",X"06C8",X"0647",X"0670",X"03F1",X"0171",X"00F8",X"0293",X"011F",X"FBA1",X"F55E",X"F215",X"F231",X"F68A",X"FFC1",X"072B",X"09D3",X"0854",X"0634",X"06A9",X"0572",X"02E0",X"00E4",X"0202",X"02B3",X"FFA5",X"F952",X"F3F8",X"F1C8",X"F2B3",X"F970",X"02B0",X"0865",X"09C4",X"0735",X"06A7",X"065E",X"0481",X"01BF",X"013D",X"02D1",X"0260",X"FDAF",X"F758",X"F348",X"F18B",X"F426",X"FCB6",X"04B6",X"0966",X"088B",X"06E3",X"06E7",X"05F1",X"0367",X"0119",X"01CA",X"02FF",X"00FC",X"FB61",X"F5EB",X"F2BC",X"F1B4",X"F71F",X"FFD3",X"071C",X"0969",X"0780",X"06D6",X"0681",X"04DA",X"01DB",X"00EB",X"028B",X"030D",X"FF9A",X"F9B9",X"F55A",X"F1F1",X"F2CE",X"F9DE",X"022D",X"0830",X"0833",X"0716",X"06DB",X"0659",X"03CF",X"0162",X"01B3",X"0351",X"025B",X"FD55",X"F82A",X"F3FC",X"F13B",X"F4F8",X"FC94",X"04FD",X"0855",X"0792",X"06F7",X"06FD",X"059F",X"02B5",X"013F",X"0283",X"0393",X"00D4",X"FB6D",X"F71F",X"F26C",X"F1EF",X"F71A",X"FFB2",X"06A8",X"07E6",X"074C",X"0739",X"06FD",X"04AA",X"01F5",X"0199",X"0330",X"0310",X"FEC0",X"FA40",X"F573",X"F1A8",X"F349",X"F9C5",X"02BE",X"0734",X"0794",X"0730",X"0767",X"0654",X"0374",X"0177",X"0216",X"03BA",X"01A8",X"FD08",X"F8C7",X"F373",X"F1A7",X"F4B0",X"FD23",X"04D6",X"0787",X"0779",X"0794",X"078F",X"0598",X"02A3",X"018B",X"030F",X"038C",X"FFB1",X"FBDA",X"F69A",X"F247",X"F1D7",X"F753",X"004A",X"061A",X"0779",X"076E",X"07C2",X"06F6",X"0439",X"01E3",X"01ED",X"03F7",X"024A",X"FEB8",X"FA7B",X"F4F2",X"F1AA",X"F306",X"FA89",X"02B1",X"06C2",X"0758",X"0792",X"07C3",X"060E",X"0313",X"013E",X"02E6",X"03CB",X"00E3",X"FDA7",X"F882",X"F3BB",X"F176",X"F54F",X"FDD4",X"04A7",X"0725",X"0780",X"0800",X"0780",X"04FD",X"01EA",X"017B",X"03AD",X"0253",X"FFBA",X"FBAC",X"F6AB",X"F23D",X"F1E9",X"F83C",X"00C5",X"0606",X"077F",X"0805",X"0848",X"06BA",X"03A3",X"00E0",X"029A",X"0372",X"01BE",X"FEC4",X"FA60",X"F552",X"F193",X"F3B0",X"FB5A",X"02C5",X"0644",X"071E",X"0801",X"07B9",X"05B2",X"020B",X"017D",X"0393",X"0308",X"0110",X"FD7E",X"F8FE",X"F3C6",X"F190",X"F61E",X"FE36",X"0416",X"063B",X"074F",X"07FE",X"0734",X"0423",X"0106",X"0292",X"037F",X"0290",X"0011",X"FC75",X"F76A",X"F28E",X"F28E",X"F8FE",X"009E",X"04E0",X"0677",X"07B3",X"07F3",X"0692",X"0263",X"01AD",X"0347",X"0369",X"01BD",X"FEC5",X"FADA",X"F553",X"F175",X"F424",X"FBAB",X"0254",X"0551",X"072E",X"080B",X"0864",X"0518",X"01DC",X"029A",X"03A5",X"0329",X"00DE",X"FDC6",X"F922",X"F361",X"F193",X"F66C",X"FE37",X"0330",X"05C5",X"0741",X"0859",X"076F",X"033A",X"0208",X"0328",X"03DE",X"026D",X"FFF5",X"FCBE",X"F733",X"F21E",X"F2BA",X"F94C",X"0045",X"0409",X"065C",X"0799",X"08AD",X"058A",X"022B",X"022C",X"0367",X"0376",X"01AE",X"FF55",X"FB54",X"F542",X"F1C8",X"F4CD",X"FC3D",X"01A8",X"0518",X"069A",X"0884",X"07E0",X"03D4",X"01EF",X"0290",X"038A",X"02B8",X"00C9",X"FE68",X"F938",X"F378",X"F1F9",X"F789",X"FE2F",X"0304",X"057D",X"0750",X"08F6",X"0646",X"02F2",X"0229",X"0360",X"03AB",X"0227",X"0058",X"FCE0",X"F6E4",X"F1D0",X"F355",X"F9BE",X"FFB9",X"03FD",X"05E7",X"089D",X"0873",X"04D5",X"023D",X"0272",X"03AE",X"0320",X"017B",X"FFBB",X"FB56",X"F4FF",X"F1EA",X"F5F2",X"FBE8",X"0187",X"0449",X"06E7",X"08F8",X"06EE",X"0351",X"01E5",X"0304",X"03C9",X"0290",X"0144",X"FEB2",X"F947",X"F306",X"F2E6",X"F7B9",X"FDFF",X"026D",X"0501",X"0830",X"0899",X"056C",X"026A",X"0229",X"039B",X"0349",X"021A",X"00B8",X"FD65",X"F6B5",X"F25D",X"F467",X"F9DB",X"FFEB",X"0303",X"063A",X"08F5",X"07AA",X"040B",X"01EF",X"02D3",X"03BA",X"02EC",X"01F0",X"0051",X"FB4A",X"F458",X"F298",X"F5C7",X"FC4E",X"00EF",X"03E7",X"079C",X"08F6",X"066E",X"02FA",X"0212",X"0376",X"0373",X"0288",X"0190",X"FF23",X"F84B",X"F300",X"F2F7",X"F7EB",X"FE0F",X"01A1",X"054F",X"08CC",X"088E",X"0531",X"0253",X"02D8",X"039D",X"031D",X"020C",X"015F",X"FCF0",X"F5F8",X"F28A",X"F468",X"FA90",X"FF62",X"02D8",X"0703",X"0927",X"0762",X"038C",X"0214",X"02FB",X"0345",X"026B",X"020C",X"00A3",X"FA83",X"F4BC",X"F2BC",X"F690",X"FC65",X"002E",X"0423",X"0804",X"08D1",X"05DA",X"027E",X"027B",X"0365",X"033F",X"0244",X"0281",X"FEDB",X"F877",X"F373",X"F3A5",X"F8DB",X"FD94",X"014D",X"05CD",X"08D2",X"081E",X"0413",X"021A",X"029B",X"0362",X"0257",X"028C",X"01B8",X"FCBA",X"F679",X"F2E9",X"F582",X"FAC8",X"FEA0",X"02C9",X"0724",X"091A",X"067C",X"02E8",X"020D",X"032C",X"02F8",X"0246",X"0310",X"0085",X"FACF",X"F4BD",X"F34C",X"F78C",X"FBEC",X"FFC5",X"044A",X"0862",X"089D",X"0509",X"0276",X"0288",X"0373",X"024A",X"02E6",X"02A4",X"FECD",X"F85A",X"F35E",X"F486",X"F909",X"FCE2",X"010C",X"05D9",X"08F8",X"0741",X"03D4",X"0223",X"0354",X"02D5",X"0279",X"036F",X"01F3",X"FD04",X"F648",X"F33D",X"F62B",X"FA31",X"FE01",X"026E",X"076A",X"08AF",X"0610",X"02B6",X"02BA",X"036B",X"027C",X"032C",X"0373",X"00DB",X"FAB3",X"F46F",X"F40B",X"F772",X"FB41",X"FF18",X"0455",X"0870",X"080E",X"048F",X"0261",X"0358",X"02C3",X"026E",X"0355",X"02CC",X"FF05",X"F7E9",X"F3B8",X"F543",X"F8DE",X"FC66",X"00DD",X"0686",X"08F6",X"0710",X"0338",X"02F1",X"0349",X"025E",X"02CA",X"037A",X"0235",X"FCB0",X"F5DD",X"F409",X"F65C",X"F9E8",X"FD6B",X"02FD",X"07BD",X"08AD",X"0523",X"02B5",X"031D",X"028B",X"023D",X"0316",X"0391",X"010E",X"FA10",X"F4E1",X"F4BF",X"F7BB",X"FABD",X"FF2E",X"04E8",X"08AA",X"07A9",X"03D7",X"0322",X"0318",X"0247",X"027A",X"036C",X"035D",X"FEB1",X"F7C1",X"F481",X"F5DA",X"F8BF",X"FBE0",X"0127",X"067A",X"08DA",X"05DE",X"0362",X"035C",X"02B2",X"0241",X"02B6",X"03E2",X"025E",X"FC14",X"F64D",X"F4BE",X"F6F7",X"F961",X"FD73",X"02E8",X"07E0",X"07D4",X"0473",X"036B",X"031B",X"0266",X"024F",X"034A",X"044D",X"0096",X"F9FB",X"F565",X"F5AE",X"F78D",X"FA4D",X"FEEF",X"04FB",X"0887",X"0663",X"03FA",X"038E",X"02E4",X"025D",X"0262",X"040E",X"036C",X"FE1F",X"F7B5",X"F530",X"F652",X"F842",X"FBB6",X"0119",X"071E",X"0836",X"0535",X"03D3",X"0338",X"02A4",X"01E9",X"02CA",X"044F",X"01DC",X"FBBA",X"F673",X"F5C9",X"F6F5",X"F956",X"FD25",X"0380",X"082B",X"06F0",X"0488",X"03A6",X"0318",X"0261",X"01F5",X"03DF",X"0411",X"0007",X"F954",X"F609",X"F60D",X"F786",X"FA09",X"FF04",X"05DE",X"080F",X"05D1",X"043C",X"037C",X"0316",X"01EA",X"02BC",X"046F",X"033E",X"FD7E",X"F7C4",X"F5DA",X"F66F",X"F838",X"FB40",X"01D5",X"076C",X"0740",X"0523",X"03C8",X"0364",X"0253",X"01A1",X"0359",X"048E",X"018D",X"FB09",X"F6FC",X"F5FA",X"F70B",X"F8CE",X"FD3C",X"047A",X"07CD",X"06A1",X"04AF",X"03BF",X"034A",X"01BF",X"0221",X"0418",X"0436",X"FF44",X"F986",X"F691",X"F689",X"F794",X"F9A3",X"FFE1",X"0634",X"0741",X"05A4",X"03DE",X"0381",X"0255",X"0178",X"02CA",X"04D7",X"02EB",X"FD3E",X"F863",X"F689",X"F702",X"F7AD",X"FB58",X"02A5",X"06DF",X"06CD",X"04AB",X"03D9",X"0341",X"01CE",X"01BF",X"03E3",X"04F0",X"0123",X"FB7A",X"F788",X"F6DB",X"F717",X"F818",X"FDFC",X"04A3",X"0723",X"05EE",X"0423",X"03BF",X"0298",X"0162",X"0239",X"04C9",X"03D4",X"FEFE",X"F9B9",X"F71F",X"F722",X"F6E0",X"F9BC",X"00CE",X"0602",X"070F",X"051B",X"042B",X"036D",X"021F",X"015C",X"0374",X"051C",X"0279",X"FD15",X"F872",X"F73C",X"F6CF",X"F6D3",X"FBFD",X"02C7",X"06BA",X"062F",X"04AA",X"0411",X"0335",X"01AE",X"0200",X"049F",X"04AA",X"00B9",X"FB1D",X"F7D3",X"F761",X"F61F",X"F81A",X"FE64",X"049E",X"06B1",X"0564",X"047E",X"03FE",X"02AC",X"014E",X"032B",X"0537",X"03B5",X"FEBA",X"F998",X"F7FA",X"F6C8",X"F603",X"FA0A",X"00E5",X"060A",X"0653",X"0508",X"0465",X"03B4",X"01BC",X"01A1",X"041C",X"0513",X"022D",X"FC79",X"F8BA",X"F7C0",X"F5DF",X"F6E3",X"FC48",X"0339",X"0660",X"05C3",X"04B3",X"0451",X"02F6",X"014A",X"02A5",X"04E5",X"04AF",X"006D",X"FAF5",X"F900",X"F723",X"F5D0",X"F843",X"FED9",X"04A8",X"0619",X"0514",X"0461",X"03E9",X"01F8",X"0169",X"0399",X"054E",X"03BD",X"FE33",X"FA4B",X"F88F",X"F64D",X"F5F7",X"FA41",X"0150",X"0585",X"05D8",X"04B8",X"0481",X"033F",X"0161",X"022E",X"0478",X"0578",X"01DF",X"FC75",X"F9FD",X"F7A1",X"F595",X"F6B8",X"FCCA",X"0337",X"05FB",X"0553",X"04B1",X"0446",X"023F",X"014B",X"0306",X"054D",X"04D4",X"FFA3",X"FBB8",X"F960",X"F6D0",X"F545",X"F869",X"FF30",X"047B",X"05A8",X"04EC",X"04E0",X"03A1",X"0198",X"01CF",X"03EE",X"0605",X"0318",X"FE21",X"FB25",X"F89F",X"F5D3",X"F5A7",X"FAAA",X"0177",X"0544",X"0532",X"04D5",X"0485",X"0286",X"0139",X"0217",X"04FD",X"0567",X"011F",X"FD2A",X"FA8B",X"F7C7",X"F542",X"F716",X"FD52",X"0375",X"057D",X"050F",X"050E",X"03E4",X"01D6",X"012B",X"0328",X"05F7",X"0401",X"FF88",X"FC2C",X"F9A6",X"F665",X"F513",X"F8D4",X"FFB3",X"0481",X"0532",X"050E",X"04DE",X"02F9",X"0161",X"016E",X"04AA",X"05C6",X"026A",X"FE6B",X"FBB8",X"F8C4",X"F594",X"F5F4",X"FB4A",X"01E7",X"04FB",X"0502",X"0537",X"0413",X"022C",X"00B7",X"0267",X"05A7",X"04CE",X"00F7",X"FD90",X"FB1A",X"F77E",X"F512",X"F758",X"FDD9",X"0370",X"04CF",X"0532",X"04F8",X"036D",X"0144",X"0094",X"03C8",X"05A5",X"036C",X"FFAD",X"FD11",X"FA0B",X"F66C",X"F565",X"F98A",X"0050",X"0421",X"04E4",X"0547",X"0469",X"02BD",X"0081",X"01B1",X"0512",X"054D",X"0214",X"FEC3",X"FC3B",X"F89B",X"F54E",X"F605",X"FBD9",X"020C",X"0435",X"053A",X"0518",X"0436",X"01D2",X"007E",X"0320",X"05B3",X"045E",X"00D2",X"FE20",X"FB32",X"F732",X"F4D2",X"F784",X"FE5E",X"02D0",X"04A1",X"053E",X"0509",X"0395",X"00CC",X"0147",X"047E",X"0594",X"02EE",X"FFD8",X"FD69",X"F9F7",X"F5FC",X"F511",X"FA18",X"0049",X"038C",X"0508",X"053B",X"04E3",X"0242",X"0052",X"023C",X"0548",X"04B5",X"01B3",X"FF22",X"FC8D",X"F893",X"F4F7",X"F654",X"FC94",X"018E",X"0438",X"0504",X"0551",X"041B",X"0120",X"00A5",X"03AF",X"0595",X"03BD",X"00D3",X"FE96",X"FB72",X"F70C",X"F47F",X"F871",X"FE69",X"028D",X"046A",X"051A",X"0544",X"02EB",X"0075",X"01A2",X"04DC",X"053D",X"02A1",X"004D",X"FDEE",X"FA43",X"F57B",X"F560",X"FAA0",X"FFF7",X"034E",X"0467",X"0560",X"04AE",X"0191",X"0031",X"02D5",X"054B",X"0434",X"01C8",X"FFBA",X"FD20",X"F88E",X"F4DE",X"F74D",X"FCA8",X"0174",X"03A7",X"04C4",X"056C",X"0382",X"0081",X"00E8",X"0424",X"0529",X"0346",X"0126",X"FF1F",X"FBDE",X"F685",X"F52F",X"F8F4",X"FE7E",X"0249",X"03D6",X"0539",X"0519",X"022B",X"0044",X"023F",X"050C",X"0490",X"027D",X"0069",X"FE68",X"F9BF",X"F54F",X"F61A",X"FAD1",X"0019",X"02DF",X"0490",X"05C6",X"044A",X"010E",X"009A",X"03A4",X"0528",X"03E5",X"01B2",X"0015",X"FD3F",X"F7B3",X"F521",X"F76B",X"FCCB",X"0108",X"032B",X"050B",X"0584",X"02E8",X"0051",X"01A8",X"0484",X"04DC",X"0325",X"0137",X"FFCC",X"FB3E",X"F654",X"F587",X"F952",X"FE98",X"01C7",X"03C3",X"0576",X"04B6",X"01A0",X"0077",X"02F7",X"04E4",X"0467",X"023A",X"0123",X"FE96",X"F93C",X"F586",X"F670",X"FB45",X"FFEB",X"0252",X"048D",X"05A5",X"03AF",X"00B9",X"0158",X"03E4",X"04F6",X"0379",X"01BA",X"00BB",X"FCAF",X"F786",X"F53F",X"F7E6",X"FD3B",X"00B9",X"031B",X"053B",X"0550",X"022F",X"0076",X"0241",X"048B",X"04A7",X"0289",X"01DE",X"FFC8",X"FAF3",X"F652",X"F5C3",X"F9DF",X"FE89",X"0151",X"03D2",X"05B3",X"043A",X"0102",X"00DE",X"0331",X"050B",X"03B8",X"025F",X"01B3",X"FE82",X"F93D",X"F59C",X"F6FF",X"FBCA",X"FF85",X"0211",X"04B5",X"0588",X"0297",X"007C",X"0176",X"041D",X"0497",X"02E6",X"0263",X"00F0",X"FCCF",X"F7B3",X"F5A9",X"F8CF",X"FD36",X"0051",X"02FE",X"0587",X"0491",X"0183",X"0097",X"0297",X"04D3",X"03ED",X"02CF",X"024C",X"FFD8",X"FAE0",X"F63A",X"F64E",X"FA49",X"FE44",X"00FA",X"040B",X"059F",X"0347",X"00EB",X"0119",X"03DB",X"04AC",X"0372",X"02F7",X"01FE",X"FE73",X"F8FD",X"F5A1",X"F782",X"FBBB",X"FF0A",X"01E6",X"050A",X"04C7",X"022A",X"0069",X"0205",X"047D",X"042E",X"0337",X"02F7",X"0133",X"FCB8",X"F745",X"F5F3",X"F919",X"FD24",X"FFDD",X"035F",X"0565",X"03E4",X"0131",X"0091",X"031E",X"046B",X"0393",X"0325",X"029B",X"0000",X"FA7E",X"F64C",X"F6EF",X"FAE9",X"FE06",X"0109",X"048F",X"0510",X"02CF",X"005E",X"016D",X"03EC",X"0404",X"0360",X"0318",X"0224",X"FE31",X"F88B",X"F5F6",X"F839",X"FC09",X"FECA",X"0297",X"052E",X"04A5",X"01A8",X"006A",X"028A",X"0417",X"03AC",X"032F",X"0305",X"014B",X"FC1E",X"F717",X"F661",X"F9C3",X"FCB4",X"000A",X"03D0",X"0560",X"0390",X"009D",X"0106",X"0351",X"03E2",X"0368",X"033A",X"0303",X"FFD6",X"FA2D",X"F655",X"F7AA",X"FAE7",X"FDA5",X"0176",X"04A7",X"0503",X"0225",X"0045",X"01F6",X"03AB",X"03B8",X"033E",X"037E",X"028E",X"FE25",X"F865",X"F66C",X"F8E3",X"FB89",X"FECB",X"02A0",X"0507",X"03EA",X"00D9",X"00AC",X"02C5",X"03D9",X"039E",X"0384",X"03D5",X"0183",X"FC15",X"F708",X"F735",X"F9B2",X"FC7D",X"0018",X"03CA",X"0513",X"02A2",X"0056",X"016B",X"032D",X"03B4",X"0346",X"03C9",X"037F",X"0011",X"F9EE",X"F6D4",X"F818",X"FA76",X"FD99",X"016E",X"04A2",X"045A",X"0145",X"0083",X"021E",X"03A5",X"0371",X"0388",X"0417",X"02F8",X"FDEE",X"F844",X"F724",X"F8B7",X"FB49",X"FEB2",X"02AC",X"04FD",X"031D",X"00B4",X"010F",X"02DC",X"03AA",X"0361",X"03D2",X"0435",X"01AC",X"FB78",X"F789",X"F78C",X"F97B",X"FC2D",X"FFF2",X"03F1",X"0497",X"01F4",X"009D",X"01C7",X"0363",X"036E",X"0372",X"040B",X"03FC",X"FF8F",X"F9BF",X"F769",X"F839",X"FA67",X"FD6C",X"01AE",X"04D3",X"03AA",X"0135",X"00B7",X"025D",X"033F",X"032B",X"036B",X"0478",X"02F1",X"FD40",X"F899",X"F7A7",X"F8DB",X"FB32",X"FEAC",X"0346",X"04BC",X"02A5",X"00B6",X"0149",X"02D3",X"0334",X"030E",X"03BE",X"0492",X"011C",X"FB59",X"F81A",X"F7FB",X"F9AB",X"FC2D",X"0091",X"044C",X"0418",X"01B5",X"009D",X"01E8",X"02E3",X"0300",X"02FF",X"048B",X"0410",X"FF26",X"FA28",X"F7F2",X"F87E",X"FA33",X"FD4F",X"0228",X"045D",X"030E",X"00D4",X"00F6",X"0239",X"0309",X"02B7",X"038F",X"050E",X"02A7",X"FD45",X"F930",X"F81A",X"F911",X"FADF",X"FF22",X"035C",X"043C",X"0209",X"00B0",X"016D",X"02BA",X"0301",X"02CD",X"0490",X"04E4",X"00CD",X"FB8E",X"F861",X"F844",X"F921",X"FBCE",X"00BA",X"0402",X"0387",X"0159",X"00EB",X"01FF",X"02FF",X"028D",X"0347",X"053E",X"03BF",X"FEF6",X"FA3D",X"F866",X"F89D",X"F9B6",X"FD9E",X"0247",X"0430",X"027C",X"0100",X"0130",X"0293",X"02EA",X"028F",X"043F",X"0550",X"0277",X"FD45",X"F963",X"F88C",X"F89B",X"FAB9",X"FF3B",X"0348",X"0384",X"01A1",X"00A6",X"019B",X"02D1",X"0250",X"02CA",X"0509",X"04B1",X"00B8",X"FBA7",X"F920",X"F885",X"F917",X"FC42",X"0112",X"03C3",X"02EB",X"0131",X"00DE",X"024F",X"02AF",X"0221",X"03C3",X"055C",X"03A4",X"FED6",X"FA93",X"F8FB",X"F87A",X"F9D9",X"FDF6",X"0279",X"038D",X"021B",X"00A8",X"013F",X"029C",X"022B",X"027E",X"049E",X"052A",X"022E",X"FCFB",X"FA02",X"F8A1",X"F892",X"FAF1",X"FFE6",X"032D",X"032E",X"0169",X"0094",X"01FD",X"0287",X"01E9",X"0347",X"0526",X"04B8",X"004C",X"FBF3",X"F99D",X"F886",X"F8FC",X"FCA8",X"0159",X"0380",X"0289",X"00B0",X"00EB",X"027B",X"0206",X"0221",X"03FD",X"0589",X"0356",X"FEAB",X"FB27",X"F930",X"F857",X"F9DF",X"FE65",X"0246",X"0341",X"01A8",X"005C",X"01B3",X"0269",X"01E8",X"02D5",X"04FE",X"057A",X"01CB",X"FD77",X"FA86",X"F8D1",X"F867",X"FB59",X"FFE9",X"02D3",X"02AD",X"00C4",X"00BD",X"0246",X"0217",X"0207",X"037B",X"05BB",X"0456",X"000B",X"FC38",X"F9F4",X"F84D",X"F902",X"FCF3",X"0126",X"0306",X"01D9",X"0069",X"0199",X"025E",X"01DC",X"0229",X"0484",X"0594",X"02D3",X"FE94",X"FB7F",X"F961",X"F855",X"FA75",X"FECB",X"024E",X"02F4",X"00E6",X"00AD",X"01E3",X"0200",X"019E",X"02DF",X"056B",X"04FF",X"016F",X"FD81",X"FAD4",X"F8AD",X"F8AD",X"FBD0",X"000A",X"02E2",X"0218",X"0073",X"013C",X"0215",X"01DD",X"01B5",X"03F2",X"05AE",X"03F0",X"FFF8",X"FCAC",X"FA0D",X"F85C",X"F992",X"FD42",X"0167",X"02EC",X"012E",X"00A0",X"0187",X"0208",X"0153",X"0249",X"04E0",X"0575",X"028E",X"FED9",X"FBE1",X"F940",X"F86B",X"FA95",X"FEB8",X"0277",X"024B",X"00CC",X"00FC",X"020C",X"01D8",X"0170",X"0356",X"0594",X"04B4",X"0130",X"FDD8",X"FAD8",X"F883",X"F8BD",X"FBB0",X"0053",X"02AD",X"0187",X"00B3",X"0174",X"022C",X"016B",X"01EA",X"0471",X"05B9",X"03A4",X"0014",X"FCDF",X"F9C5",X"F84A",X"F974",X"FD42",X"0198",X"0245",X"0102",X"00C3",X"01E2",X"01D3",X"013D",X"02AE",X"0550",X"0562",X"0286",X"FF42",X"FBF8",X"F91B",X"F874",X"FA6B",X"FF28",X"021E",X"01B2",X"008D",X"0114",X"01EE",X"014D",X"015E",X"03BA",X"05B3",X"0469",X"016A",X"FE25",X"FAB5",X"F8B4",X"F8B7",X"FC17",X"00AF",X"0252",X"0148",X"00B2",X"01AE",X"01CD",X"010A",X"0202",X"04D9",X"0588",X"0367",X"0078",X"FCEC",X"F9E9",X"F85A",X"F969",X"FDE2",X"0182",X"01DD",X"00AC",X"00F3",X"01E2",X"0170",X"0101",X"0316",X"057B",X"0503",X"028E",X"FF52",X"FBB2",X"F93A",X"F827",X"FACD",X"FF69",X"01E7",X"0148",X"0095",X"0179",X"01E5",X"00FA",X"0199",X"0451",X"05B1",X"043C",X"01B1",X"FE04",X"FAE3",X"F888",X"F8CB",X"FC91",X"00C9",X"01EC",X"00C9",X"00C4",X"01B3",X"0158",X"00A0",X"0240",X"04DF",X"050F",X"036C",X"0068",X"FCF7",X"FA11",X"F84B",X"FA0D",X"FE7E",X"01BF",X"018E",X"00A0",X"0136",X"01B4",X"00C4",X"00DA",X"0365",X"0521",X"04AE",X"029F",X"FF43",X"FC16",X"F91D",X"F873",X"FB61",X"FFE5",X"01D4",X"0110",X"00BC",X"01A6",X"016D",X"0078",X"01A7",X"043D",X"0520",X"0463",X"0198",X"FE4C",X"FAF9",X"F873",X"F900",X"FCF7",X"00D3",X"0173",X"0089",X"00F9",X"01B9",X"00E9",X"0080",X"02BE",X"04B6",X"054B",X"03A3",X"00A1",X"FD73",X"FA08",X"F847",X"FA3A",X"FE9E",X"0142",X"00F2",X"0089",X"0151",X"0172",X"0056",X"013C",X"0380",X"0501",X"04E5",X"029B",X"FFA6",X"FC4F",X"F93E",X"F89B",X"FBBD",X"FFD6",X"013C",X"0081",X"00C2",X"01B0",X"00F4",X"004E",X"021E",X"041C",X"054C",X"0439",X"01A3",X"FE8C",X"FB0B",X"F871",X"F945",X"FD56",X"00B5",X"00FD",X"008C",X"0163",X"01B4",X"0069",X"00FA",X"02D1",X"04B7",X"0522",X"0360",X"00BC",X"FD6D",X"F9DC",X"F83E",X"FA7A",X"FEB2",X"00C8",X"007C",X"0097",X"01B3",X"0106",X"006B",X"0198",X"0394",X"053F",X"04CF",X"02C5",X"FFE7",X"FC5A",X"F906",X"F8AB",X"FC13",X"FFD0",X"00B7",X"002E",X"010E",X"0177",X"005E",X"0084",X"0200",X"0437",X"0536",X"0443",X"01E7",X"FEE5",X"FB22",X"F893",X"F9AF",X"FDC1",X"0085",X"007C",X"0081",X"0196",X"00F8",X"0038",X"00BE",X"02A4",X"04A8",X"0508",X"0382",X"0107",X"FDAC",X"F9E1",X"F86B",X"FB24",X"FF10",X"009E",X"0029",X"0111",X"0165",X"0096",X"0050",X"0158",X"0393",X"051B",X"04BC",X"02DD",X"001B",X"FC51",X"F8D5",X"F8F8",X"FC6D",X"FFBF",X"001A",X"0058",X"015E",X"0110",X"0068",X"0088",X"0225",X"0458",X"053E",X"0440",X"0219",X"FF01",X"FAFB",X"F894",X"FA1D",X"FE0F",X"0016",X"FFFD",X"00C9",X"012B",X"0091",X"0000",X"00C0",X"02CF",X"04BE",X"04FE",X"03AD",X"015E",X"FDD2",X"F9DB",X"F8BF",X"FB93",X"FF18",X"FFD8",X"0042",X"0116",X"0113",X"0069",X"0034",X"016A",X"03AE",X"04FC",X"049A",X"02DA",X"0042",X"FC2B",X"F8F7",X"F94D",X"FD20",X"FF72",X"FFCE",X"00B3",X"0147",X"0100",X"005A",X"008B",X"0242",X"0456",X"0516",X"0414",X"023B",X"FEFD",X"FACB",X"F881",X"FA94",X"FE3A",X"FF5C",X"0007",X"00DD",X"0115",X"0098",X"0034",X"00F6",X"0301",X"04B7",X"04C3",X"038F",X"0152",X"FD8F",X"F9B1",X"F8F1",X"FC42",X"FED0",X"FF93",X"0062",X"0117",X"0100",X"0064",X"0038",X"0199",X"03AD",X"04EB",X"046A",X"0303",X"0045",X"FC2F",X"F8DC",X"FA22",X"FD69",X"FF13",X"FFE2",X"00AE",X"00E6",X"00AF",X"0010",X"0068",X"0233",X"044A",X"04C4",X"0415",X"0241",X"FF04",X"FAA1",X"F8E0",X"FB6C",X"FE12",X"FF51",X"0035",X"00CB",X"00EE",X"0074",X"002D",X"010A",X"0333",X"04BB",X"04CC",X"03BC",X"017F",X"FD84",X"F963",X"F992",X"FC52",X"FE59",X"FF78",X"004E",X"00B6",X"00B0",X"0017",X"0029",X"01B1",X"03E8",X"04EE",X"04A3",X"0337",X"008C",X"FBBE",X"F90F",X"FA93",X"FD28",X"FEB8",X"FFC5",X"0069",X"00CB",X"007A",X"0009",X"007E",X"029F",X"0464",X"04F4",X"0446",X"02BE",X"FF03",X"FA50",X"F967",X"FBA1",X"FDC7",X"FF2F",X"000B",X"00A8",X"00A5",X"0037",X"FFE7",X"0113",X"0339",X"04BD",X"04BF",X"03DD",X"01CB",X"FD08",X"F96D",X"F9FD",X"FC52",X"FE34",X"FF66",X"0038",X"00B5",X"00B5",X"0030",X"0046",X"01EF",X"03E6",X"04DD",X"046F",X"0399",X"0049",X"FB5D",X"F970",X"FAED",X"FD0B",X"FEB5",X"FFCD",X"0086",X"00C8",X"0071",X"FFDF",X"009E",X"027E",X"0459",X"04A3",X"0462",X"02E8",X"FE7D",X"FA4B",X"F9DE",X"FB9C",X"FDA3",X"FF11",X"001A",X"0086",X"00A6",X"0002",X"FFE5",X"011C",X"0354",X"048B",X"0493",X"0461",X"01C2",X"FCB8",X"F9FC",X"FA81",X"FC79",X"FE2E",X"FF87",X"003E",X"00A6",X"006C",X"FFC0",X"0014",X"01D1",X"03E6",X"0465",X"049E",X"03E5",X"FFEB",X"FB60",X"F9E7",X"FB28",X"FD1A",X"FEC6",X"FFE6",X"0082",X"00C1",X"001A",X"FFBC",X"0075",X"02B0",X"041B",X"0460",X"04D5",X"02E4",X"FE30",X"FAB4",X"FA55",X"FBEE",X"FDBB",X"FF47",X"0000",X"008B",X"005A",X"FFC4",X"FF9B",X"012E",X"0367",X"0432",X"04B5",X"04A7",X"0142",X"FCAA",X"FA41",X"FAD5",X"FC89",X"FE5E",X"FF8A",X"0049",X"008F",X"0026",X"FF78",X"FFDE",X"0219",X"03AC",X"0441",X"0525",X"03F7",X"FFA8",X"FBA9",X"FA71",X"FB5B",X"FD3B",X"FED2",X"FFC5",X"0063",X"005F",X"FFE5",X"FF55",X"0099",X"02D7",X"03CF",X"04C5",X"052E",X"0294",X"FDF7",X"FACD",X"FA7E",X"FBD8",X"FDC9",X"FF19",X"0013",X"0072",X"005D",X"FF87",X"FF89",X"0190",X"0345",X"0401",X"0543",X"04B4",X"010C",X"FCAA",X"FA94",X"FADA",X"FC99",X"FE49",X"FF88",X"002D",X"0083",X"0014",X"FF39",X"0015",X"024F",X"0350",X"0476",X"055F",X"03A8",X"FF57",X"FBBC",X"FA7F",X"FB5E",X"FD30",X"FEB3",X"FFC5",X"0053",X"0088",X"FFA5",X"FF45",X"0112",X"02B8",X"0396",X"0505",X"0538",X"0241",X"FDEA",X"FB11",X"FA97",X"FC05",X"FDBF",X"FF34",X"FFF3",X"007C",X"0045",X"FF39",X"FFBE",X"01BB",X"02DA",X"0414",X"056A",X"047B",X"00B3",X"FCD2",X"FAA3",X"FB0D",X"FC9F",X"FE5F",X"FF7F",X"0022",X"009C",X"FFD3",X"FF0B",X"007B",X"0204",X"031D",X"04AC",X"0598",X"0370",X"FF6E",X"FBF6",X"FABD",X"FB80",X"FD31",X"FED7",X"FFB1",X"006B",X"007D",X"FF39",X"FF6D",X"010A",X"022E",X"0356",X"051E",X"050F",X"0212",X"FE19",X"FB54",X"FAE5",X"FC07",X"FDDE",X"FF25",X"FFE8",X"00C1",X"FFFF",X"FF06",X"0011",X"0194",X"028A",X"0423",X"059B",X"0448",X"00C9",X"FCF9",X"FB06",X"FB20",X"FC8E",X"FE3F",X"FF2C",X"003E",X"00A7",X"FF5F",X"FF5F",X"00C0",X"01D7",X"0311",X"04FB",X"0564",X"033A",X"FF4F",X"FC21",X"FADD",X"FB89",X"FD42",X"FE90",X"FF86",X"00A2",X"001A",X"FF20",X"FFBA",X"010F",X"01F3",X"03AD",X"055D",X"04F0",X"0209",X"FE32",X"FB9F",X"FB0E",X"FC42",X"FDF0",X"FED6",X"001F",X"009D",X"FF77",X"FF22",X"003E",X"013C",X"025A",X"0471",X"0578",X"042A",X"00B4",X"FD22",X"FB2D",X"FB50",X"FCF5",X"FE28",X"FF2F",X"0094",X"001C",X"FF11",X"FF7C",X"00B2",X"016A",X"031E",X"0502",X"0562",X"0318",X"FF64",X"FC46",X"FAF7",X"FBD8",X"FD79",X"FE54",X"FFCB",X"009B",X"FFAC",X"FF04",X"0000",X"00D5",X"01E7",X"03D6",X"0560",X"04D0",X"01E6",X"FE4D",X"FBAD",X"FB29",X"FC9D",X"FDAA",X"FECA",X"004A",X"0038",X"FEFB",X"FF3E",X"0032",X"010C",X"0288",X"0494",X"0589",X"0413",X"00BB",X"FD53",X"FB38",X"FBB2",X"FD0E",X"FDE9",X"FF6F",X"007F",X"FFAB",X"FEFC",X"FFB5",X"006F",X"016D",X"0339",X"0517",X"054B",X"0309",X"FF93",X"FC66",X"FB34",X"FC48",X"FD2C",X"FE4C",X"FFEA",X"0045",X"FF1C",X"FF2B",X"FFF1",X"00B6",X"01F4",X"03F5",X"0571",X"04B6",X"01F7",X"FE7F",X"FBA8",X"FBA4",X"FCA7",X"FD7B",X"FEE8",X"0058",X"FFC2",X"FF00",X"FF68",X"0027",X"00F2",X"029C",X"04AB",X"057A",X"03E7",X"00F7",X"FD42",X"FB8D",X"FC22",X"FCEE",X"FDDD",X"FF95",X"0026",X"FF34",X"FEF8",X"FF90",X"003E",X"0156",X"0355",X"052C",X"050F",X"0327",X"FFAB",X"FC57",X"FBB4",X"FC6C",X"FD20",X"FE88",X"0019",X"FFBF",X"FEF4",X"FF27",X"FFDF",X"0090",X"0208",X"0437",X"0575",X"04A4",X"0227",X"FE4B",X"FBE5",X"FBF1",X"FC9C",X"FD61",X"FF54",X"001C",X"FF58",X"FEF0",X"FF69",X"FFF8",X"00D0",X"02AE",X"04D5",X"053A",X"0417",X"00D3",X"FD2D",X"FBBD",X"FC38",X"FC99",X"FE02",X"FFC4",X"FFD9",X"FF17",X"FF1B",X"FFA2",X"0032",X"015D",X"039E",X"052C",X"052D",X"0353",X"FF70",X"FC78",X"FC01",X"FC3B",X"FCCB",X"FEC6",X"0003",X"FF90",X"FF00",X"FF3E",X"FFC2",X"0053",X"0206",X"043A",X"052B",X"04D7",X"020B",X"FE28",X"FC30",X"FC2F",X"FC31",X"FD8D",X"FF70",X"FFEB",X"FF3A",X"FF05",X"FF66",X"FFE1",X"00CB",X"02F5",X"0497",X"0555",X"042F",X"00AC",X"FD3C",X"FC49",X"FC17",X"FC84",X"FE5D",X"FFD1",X"FF97",X"FF07",X"FF1D",X"FF9C",X"FFED",X"017E",X"038E",X"04F7",X"053D",X"0321",X"FF30",X"FCCB",X"FC2D",X"FC00",X"FD1E",X"FF1B",X"FFD6",X"FF61",X"FEFB",X"FF65",X"FF89",X"004A",X"0241",X"0402",X"053E",X"04E8",X"01C5",X"FE2D",X"FCB5",X"FC18",X"FC4A",X"FDF6",X"FF8B",X"FFA7",X"FEFE",X"FEFA",X"FF4B",X"FF82",X"00F7",X"02DC",X"0476",X"0565",X"041A",X"0054",X"FD99",X"FC8C",X"FC1E",X"FCE3",X"FEC1",X"FFBE",X"FF6F",X"FEC5",X"FF14",X"FF1A",X"FFDC",X"019D",X"0360",X"04D8",X"0571",X"02D9",X"FF27",X"FD46",X"FC5E",X"FC2A",X"FD87",X"FF3C",X"FFCB",X"FF16",X"FEFB",X"FF18",X"FF39",X"0073",X"023C",X"03ED",X"0571",X"04D0",X"0150",X"FE50",X"FCD9",X"FBFF",X"FC78",X"FE2E",X"FF98",X"FF7C",X"FEFE",X"FF0F",X"FEF8",X"FF96",X"0123",X"02C3",X"0490",X"05C1",X"03C9",X"003F",X"FDE5",X"FC7E",X"FBF0",X"FD00",X"FEC0",X"FFA0",X"FF1E",X"FF10",X"FEFE",X"FEF7",X"0014",X"01A8",X"033F",X"054C",X"056F",X"0286",X"FF51",X"FD74",X"FC24",X"FC3D",X"FDA5",X"FF5C",X"FF6B",X"FF0B",X"FF04",X"FEDA",X"FF3E",X"00A4",X"01FD",X"03F5",X"05AF",X"049A",X"0141",X"FEB2",X"FCDD",X"FBFE",X"FC90",X"FE73",X"FF7E",X"FF56",X"FF30",X"FEFE",X"FEDD",X"FFBB",X"0116",X"0283",X"04CF",X"05A9",X"0361",X"0052",X"FE01",X"FC6A",X"FC00",X"FD35",X"FF08",X"FF5D",X"FF36",X"FF10",X"FEC9",X"FF07",X"0038",X"014D",X"0357",X"0577",X"0526",X"0264",X"FFA1",X"FD70",X"FC28",X"FC2E",X"FDFF",X"FF4E",X"FF5F",X"FF37",X"FEF7",X"FE92",X"FF5F",X"0071",X"01B8",X"0427",X"05CB",X"043E",X"017A",X"FED4",X"FCEE",X"FBE8",X"FCD8",X"FEA5",X"FF59",X"FF53",X"FF2F",X"FE97",X"FEBB",X"FFDA",X"00C3",X"0280",X"051D",X"056B",X"035C",X"008C",X"FE2A",X"FC78",X"FC18",X"FD91",X"FF07",X"FF46",X"FF4D",X"FEF1",X"FE6E",X"FF17",X"000A",X"011D",X"037F",X"0585",X"04E9",X"0274",X"FFB9",X"FD7D",X"FBF4",X"FC6E",X"FE35",X"FF24",X"FF4C",X"FF51",X"FE9A",X"FE9C",X"FF7E",X"002F",X"01BB",X"048B",X"0591",X"043B",X"018E",X"FF19",X"FCDF",X"FBFE",X"FD2D",X"FEB2",X"FF23",X"FF76",X"FEFC",X"FE5C",X"FEE2",X"FFC8",X"0072",X"02D1",X"052D",X"0558",X"0349",X"00B1",X"FE48",X"FC3D",X"FC31",X"FDC2",X"FEB7",X"FF3B",X"FF5D",X"FE9E",X"FE71",X"FF64",X"FFC5",X"012B",X"03C4",X"0577",X"04D4",X"027A",X"FFFD",X"FD6F",X"FC06",X"FCD1",X"FE42",X"FEE7",X"FF74",X"FF0B",X"FE44",X"FEC8",X"FF6F",X"FFEC",X"0203",X"0477",X"0576",X"0407",X"01CC",X"FF2B",X"FCC0",X"FC38",X"FD85",X"FE7C",X"FF44",X"FF81",X"FE9F",X"FE4F",X"FF1A",X"FF59",X"0066",X"02C0",X"0514",X"050D",X"0353",X"0105",X"FE3C",X"FC5A",X"FCBF",X"FDF0",X"FED3",X"FF8F",X"FF40",X"FE3F",X"FEAB",X"FF2B",X"FF7E",X"0108",X"03B1",X"053A",X"0476",X"0298",X"001C",X"FD52",X"FC4D",X"FD34",X"FE32",X"FF1B",X"FFB3",X"FECB",X"FE4D",X"FEFA",X"FF26",X"FFD0",X"01EF",X"048A",X"0518",X"03EF",X"01EE",X"FF1B",X"FCB6",X"FC97",X"FD81",X"FE79",X"FF80",X"FF62",X"FE57",X"FEA6",X"FF12",X"FF3D",X"0052",X"02FD",X"04F0",X"04BC",X"034E",X"010A",X"FDFF",X"FC81",X"FCFC",X"FDDD",X"FEF1",X"FFCA",X"FEDF",X"FE68",X"FED5",X"FF10",X"FF4B",X"012A",X"03CD",X"04F3",X"044C",X"02BA",X"FFE0",X"FD3B",X"FCA7",X"FD4F",X"FE1E",X"FF88",X"FF90",X"FE92",X"FE93",X"FF15",X"FF14",X"FFC7",X"021F",X"045A",X"04BF",X"03E0",X"01E1",X"FEC5",X"FCF5",X"FD05",X"FD7C",X"FEA9",X"FFC0",X"FEFE",X"FE7A",X"FEBC",X"FF08",X"FF08",X"0068",X"0305",X"04A1",X"048A",X"0386",X"00D8",X"FDF3",X"FCEC",X"FD1D",X"FDBD",X"FF49",X"FF77",X"FEAB",X"FE6E",X"FEF3",X"FEE0",X"FF41",X"014D",X"03C6",X"0498",X"0463",X"02C4",X"FFC3",X"FD87",X"FD27",X"FD30",X"FE7F",X"FFA4",X"FF32",X"FE54",X"FE96",X"FEE0",X"FEC1",X"FFC0",X"0242",X"0415",X"049A",X"041D",X"01CF",X"FEB7",X"FD71",X"FD17",X"FD90",X"FF1E",X"FF93",X"FED8",X"FE61",X"FECF",X"FECC",X"FEDB",X"0093",X"0309",X"044B",X"049F",X"0387",X"0090",X"FE19",X"FD47",X"FCF8",X"FE15",X"FF59",X"FF51",X"FE6F",X"FE8F",X"FEE6",X"FEC3",X"FF4F",X"0196",X"0385",X"048A",X"0495",X"02B0",X"FF8B",X"FDF0",X"FD0D",X"FD35",X"FEA0",X"FF81",X"FED3",X"FE4B",X"FEAA",X"FED0",X"FE9B",X"0019",X"025B",X"03EF",X"04BF",X"044C",X"0191",X"FF0F",X"FDAE",X"FCF3",X"FDC4",X"FF2F",X"FF46",X"FE5E",X"FE4F",X"FEAD",X"FE77",X"FEDB",X"00D4",X"02E6",X"042D",X"04E9",X"037D",X"0089",X"FE9E",X"FD3A",X"FD1E",X"FE6B",X"FF7E",X"FF01",X"FE61",X"FE97",X"FEBC",X"FE64",X"FF86",X"01A5",X"034C",X"0496",X"04BC",X"0248",X"FFCE",X"FDF6",X"FCFF",X"FD74",X"FEFC",X"FF68",X"FE98",X"FE3B",X"FEAE",X"FE5D",X"FE93",X"0059",X"025A",X"03C5",X"0522",X"040A",X"0161",X"FF30",X"FD92",X"FCEC",X"FE07",X"FF4B",X"FF19",X"FE4E",X"FE7C",X"FE9D",X"FE3B",X"FF06",X"010A",X"0299",X"0460",X"04FC",X"0318",X"00AB",X"FEAD",X"FD44",X"FD63",X"FECC",X"FF7E",X"FECF",X"FE46",X"FE92",X"FE49",X"FE2E",X"FF98",X"0169",X"0306",X"04EB",X"0465",X"0244",X"0007",X"FE26",X"FD21",X"FDED",X"FF4D",X"FF66",X"FE8B",X"FE88",X"FE8C",X"FE0C",X"FE83",X"0044",X"01C2",X"03EF",X"04F8",X"03AD",X"0179",X"FF59",X"FD87",X"FD39",X"FE6D",X"FF89",X"FEFA",X"FE87",X"FEA5",X"FE67",X"FE17",X"FF5A",X"00BD",X"0283",X"048D",X"04BC",X"02FF",X"00C7",X"FE9E",X"FD23",X"FD79",X"FF01",X"FF4B",X"FE94",X"FE61",X"FE80",X"FDFB",X"FE6F",X"FFCC",X"011C",X"0370",X"04FB",X"0461",X"0250",X"0033",X"FE17",X"FD27",X"FE23",X"FF64",X"FF0E",X"FE75",X"FE8F",X"FE42",X"FDD1",X"FEF0",X"0004",X"01D5",X"0419",X"04E1",X"03A2",X"019F",X"FF58",X"FD86",X"FD57",X"FED4",X"FF6B",X"FECC",X"FE96",X"FEB0",X"FDE2",X"FE4B",X"FF41",X"0069",X"0299",X"0498",X"0482",X"0305",X"00D5",X"FE90",X"FD18",X"FDDF",X"FF39",X"FF3E",X"FEA7",X"FECF",X"FE55",X"FDF7",X"FEBB",X"FF88",X"0112",X"0382",X"04C7",X"0418",X"0258",X"0025",X"FDDD",X"FD2E",X"FE64",X"FF4D",X"FEDB",X"FEAC",X"FEB1",X"FDE3",X"FE2D",X"FEE8",X"FFD1",X"01DF",X"042E",X"04BB",X"03AA",X"01C3",X"FF64",X"FD72",X"FDBA",X"FF06",X"FF3E",X"FEAC",X"FEE6",X"FE44",X"FDDF",X"FE6C",X"FF0A",X"004B",X"02C8",X"0482",X"0471",X"030A",X"0108",X"FE64",X"FD49",X"FE34",X"FF4C",X"FEDA",X"FEEF",X"FEB8",X"FDF9",X"FE1C",X"FEAA",X"FF40",X"0124",X"0370",X"0496",X"03FD",X"0283",X"0015",X"FDC0",X"FD81",X"FECB",X"FF23",X"FEE1",X"FF12",X"FE73",X"FE01",X"FE5F",X"FEC1",X"FFB9",X"01F8",X"040B",X"0483",X"039A",X"01CD",X"FF23",X"FD73",X"FDF6",X"FF17",X"FEE9",X"FF03",X"FED6",X"FE14",X"FE08",X"FE6B",X"FEC6",X"005F",X"02C1",X"0462",X"0454",X"034D",X"0102",X"FE62",X"FD72",X"FEA6",X"FF05",X"FEF3",X"FF0D",X"FE72",X"FDEE",X"FE42",X"FE69",X"FF2F",X"012A",X"037D",X"045E",X"042A",X"02A8",X"0000",X"FDBB",X"FDF5",X"FEF6",X"FEE9",X"FF24",X"FEED",X"FE22",X"FE17",X"FE57",X"FE7D",X"FFA1",X"0208",X"03E5",X"0464",X"03CE",X"01D5",X"FEE9",X"FD8A",X"FE77",X"FEE1",X"FF13",X"FF45",X"FE99",X"FE00",X"FE30",X"FE43",X"FEB2",X"006B",X"02DD",X"0428",X"0479",X"0370",X"00ED",X"FE1D",X"FDF1",X"FEAD",X"FED8",X"FF26",X"FF0F",X"FE39",X"FE09",X"FE29",X"FE43",X"FF02",X"0155",X"034F",X"0452",X"0426",X"02C0",X"FF9E",X"FDE1",X"FE61",X"FEC4",X"FF08",X"FF74",X"FEB5",X"FE19",X"FE1B",X"FE39",X"FE4A",X"FFC4",X"020D",X"03BB",X"0451",X"0412",X"01CA",X"FEC6",X"FE15",X"FE99",X"FEB5",X"FF43",X"FF2F",X"FE66",X"FE11",X"FE39",X"FE13",X"FE94",X"008D",X"02B4",X"040A",X"046F",X"039D",X"007E",X"FE55",X"FE51",X"FE94",X"FEEF",X"FF59",X"FEC1",X"FE22",X"FE0C",X"FE2F",X"FDFB",X"FF1C",X"013D",X"0336",X"042D",X"0495",X"02AA",X"FF85",X"FE68",X"FEA0",X"FEAE",X"FF53",X"FF46",X"FE92",X"FE05",X"FE3D",X"FDFB",X"FE35",X"FFBC",X"01FE",X"0363",X"046B",X"0419",X"0152",X"FED1",X"FE7E",X"FE77",X"FEDD",X"FF67",X"FF15",X"FE4C",X"FE3B",X"FE3E",X"FE06",X"FEB5",X"00B7",X"0292",X"03D4",X"04C2",X"0344",X"0022",X"FE9E",X"FE65",X"FE82",X"FF1A",X"FF59",X"FEB4",X"FE2B",X"FE49",X"FE0E",X"FE19",X"FF4A",X"0168",X"02E4",X"045C",X"049C",X"0210",X"FF77",X"FEA6",X"FE62",X"FED3",X"FF5E",X"FF36",X"FE54",X"FE41",X"FE2A",X"FDF0",X"FE42",X"001E",X"01DC",X"0347",X"04C6",X"03FB",X"00F8",X"FF2F",X"FE81",X"FE82",X"FF16",X"FF83",X"FED3",X"FE3D",X"FE3A",X"FE17",X"FDD3",X"FEDB",X"00BA",X"022F",X"03F7",X"04D3",X"02C1",X"0027",X"FEEF",X"FE74",X"FEA8",X"FF76",X"FF5C",X"FE80",X"FE3E",X"FE2D",X"FDE6",X"FE00",X"FF9A",X"012E",X"02B4",X"04A8",X"047A",X"01D4",X"FFC0",X"FEAD",X"FE79",X"FEFD",X"FF96",X"FF00",X"FE5E",X"FE3A",X"FE2B",X"FDAA",X"FE7F",X"0029",X"0192",X"0387",X"050D",X"037B",X"010F",X"FF4D",X"FE80",X"FE7E",X"FF59",X"FF65",X"FEA4",X"FE31",X"FE4C",X"FDDA",X"FDCA",X"FF26",X"009A",X"0217",X"046E",X"04AB",X"0293",X"0058",X"FF0B",X"FE73",X"FEF5",X"FF8F",X"FF2F",X"FE74",X"FE49",X"FE3D",X"FDA7",X"FE30",X"FF9D",X"00C6",X"02E3",X"04CA",X"0405",X"01BF",X"FFE0",X"FEBB",X"FE7B",X"FF4D",X"FF77",X"FECD",X"FE3A",X"FE59",X"FDEF",X"FDBB",X"FEDF",X"FFEB",X"015D",X"03DF",X"04CE",X"034D",X"0112",X"FF8F",X"FE81",X"FEE3",X"FF82",X"FF56",X"FE70",X"FE50",X"FE35",X"FDA3",X"FDF7",X"FF36",X"0006",X"0235",X"047D",X"047B",X"027F",X"00A1",X"FF17",X"FE9B",X"FF33",X"FF9B",X"FEF4",X"FE57",X"FE61",X"FDEE",X"FD84",X"FE8B",X"FF55",X"00AC",X"033B",X"04CE",X"03C6",X"01C3",X"FFF6",X"FEB2",X"FEC1",X"FF7B",X"FF86",X"FEAF",X"FE74",X"FE5B",X"FD90",X"FDE4",X"FEEA",X"FF96",X"0189",X"0409",X"04A6",X"030C",X"0124",X"FF59",X"FE96",X"FF07",X"FFB5",X"FF31",X"FE91",X"FE92",X"FE0E",X"FD7A",X"FE5F",X"FEDE",X"0001",X"0277",X"0488",X"041B",X"027C",X"0084",X"FEF2",X"FEA5",X"FF67",X"FFA6",X"FEE0",X"FE8D",X"FE81",X"FD87",X"FDB6",X"FE75",X"FF09",X"00C6",X"0396",X"04AE",X"03B3",X"01ED",X"FFE5",X"FEA9",X"FEF6",X"FFBE",X"FF5E",X"FE9A",X"FEA8",X"FDF0",X"FD60",X"FE04",X"FE94",X"FF5B",X"01CA",X"0434",X"0473",X"032A",X"0129",X"FF63",X"FEA6",X"FF61",X"FFC3",X"FEF5",X"FEBA",X"FE95",X"FDA1",X"FDBE",X"FE4D",X"FE9F",X"FFF7",X"02D4",X"0460",X"0408",X"027E",X"006E",X"FED8",X"FED4",X"FFB6",X"FF82",X"FEC8",X"FEEC",X"FE1C",X"FD8C",X"FDFF",X"FE6C",X"FED7",X"00FF",X"0389",X"047B",X"0391",X"01C3",X"FFAD",X"FE9E",X"FF37",X"FFDE",X"FF19",X"FEFD",X"FEB3",X"FDC3",X"FDA6",X"FE2C",X"FE48",X"FF5A",X"0202",X"0419",X"0457",X"0322",X"0112",X"FF34",X"FED4",X"FFBF",X"FFAD",X"FF10",X"FF11",X"FE3E",X"FD8D",X"FDDE",X"FE2A",X"FE3C",X"0028",X"02BF",X"043A",X"03F1",X"0270",X"004D",X"FED8",X"FF41",X"FFF6",X"FF53",X"FF47",X"FEEE",X"FDF9",X"FDA4",X"FE29",X"FDFB",X"FECE",X"011C",X"0366",X"0432",X"0387",X"01B6",X"FFA0",X"FECD",X"FFBC",X"FFAA",X"FF44",X"FF3C",X"FE83",X"FDA4",X"FDF3",X"FE1E",X"FDFA",X"FF6A",X"01FB",X"03D6",X"042E",X"031C",X"010C",X"FF0F",X"FF3F",X"FFCC",X"FF62",X"FF51",X"FF0B",X"FE03",X"FDB4",X"FE1B",X"FDD4",X"FE39",X"0038",X"02B7",X"0417",X"0402",X"0296",X"0041",X"FF12",X"FFBB",X"FF9C",X"FF64",X"FF6A",X"FEB5",X"FDB8",X"FDF3",X"FE02",X"FDB8",X"FEAD",X"0116",X"033D",X"041E",X"0399",X"01B5",X"FF66",X"FF56",X"FFB9",X"FF75",X"FF8A",X"FF68",X"FE53",X"FDF3",X"FE3D",X"FDF4",X"FDF0",X"FF7F",X"01E6",X"03A2",X"0406",X"0325",X"00AC",X"FF44",X"FF8E",X"FF9B",X"FF6A",X"FF91",X"FEEC",X"FDF8",X"FE17",X"FE31",X"FDC8",X"FE55",X"005F",X"02C2",X"03EE",X"0413",X"0258",X"FFE2",X"FF4A",X"FFA2",X"FF6F",X"FF76",X"FF6C",X"FE6A",X"FDEC",X"FE2E",X"FDE9",X"FDAA",X"FEE0",X"0138",X"032D",X"042E",X"03D0",X"015A",X"FFB1",X"FFA3",X"FFA8",X"FF76",X"FFC1",X"FF18",X"FE14",X"FE08",X"FE15",X"FDA1",X"FDD5",X"FF8A",X"01EA",X"038A",X"0462",X"02F5",X"0072",X"FF8E",X"FFB0",X"FF80",X"FFB1",X"FFBC",X"FEA9",X"FE00",X"FE33",X"FDE9",X"FD8C",X"FE44",X"0076",X"026E",X"0404",X"0425",X"01FC",X"0000",X"FFC4",X"FFA9",X"FF86",X"FFE0",X"FF4F",X"FE3D",X"FE0B",X"FE1F",X"FDB4",X"FD98",X"FF08",X"0124",X"0301",X"046F",X"0376",X"0118",X"FFF1",X"FFCA",X"FF8D",X"FFC1",X"FFD6",X"FEDB",X"FE14",X"FE22",X"FE00",X"FD85",X"FDE1",X"FFD2",X"01A1",X"03B9",X"0465",X"029B",X"007C",X"FFFF",X"FFA9",X"FF95",X"FFF8",X"FF94",X"FE6A",X"FE28",X"FE2B",X"FDCC",X"FD53",X"FE8C",X"004F",X"0246",X"0435",X"03DE",X"0193",X"003E",X"FFEC",X"FF97",X"FFD4",X"000D",X"FF12",X"FE3B",X"FE35",X"FE29",X"FD70",X"FD9D",X"FF29",X"00DF",X"0329",X"0482",X"032A",X"0113",X"003D",X"FFB9",X"FF92",X"0006",X"FFB1",X"FE9F",X"FE2C",X"FE57",X"FDF8",X"FD5A",X"FE34",X"FF98",X"018A",X"03D6",X"0437",X"0235",X"00B3",X"001A",X"FF93",X"FFD0",X"0033",X"FF50",X"FE62",X"FE39",X"FE46",X"FD79",X"FD87",X"FE9E",X"001E",X"0273",X"0465",X"0377",X"018F",X"0087",X"FFE7",X"FF99",X"002C",X"FFEE",X"FEEC",X"FE2D",X"FE6B",X"FDF4",X"FD5C",X"FDE1",X"FF04",X"00C5",X"036C",X"0448",X"02B1",X"0129",X"004F",X"FF9A",X"FFD4",X"002F",X"FF98",X"FE85",X"FE4C",X"FE5B",X"FD94",X"FD87",X"FE47",X"FF87",X"01D2",X"0421",X"03D7",X"021D",X"00E6",X"0001",X"FF98",X"0011",X"0012",X"FF2D",X"FE44",X"FE71",X"FDF9",X"FD6C",X"FDBA",X"FE88",X"000F",X"02D9",X"043C",X"032D",X"019B",X"0098",X"FFA9",X"FFDF",X"0040",X"FFEB",X"FEB6",X"FE65",X"FE5A",X"FDAA",X"FD70",X"FE04",X"FECE",X"0109",X"03A0",X"03FE",X"0278",X"0166",X"002B",X"FFBE",X"0026",X"0065",X"FF71",X"FE81",X"FE8B",X"FE22",X"FD76",X"FDA6",X"FE26",X"FF5A",X"0213",X"0406",X"0360",X"0210",X"00D2",X"FFDA",X"FFC5",X"0057",X"0038",X"FEF4",X"FE8E",X"FE7D",X"FDCA",X"FD83",X"FDCA",X"FE40",X"0038",X"030B",X"03F1",X"02ED",X"01C0",X"0065",X"FFC2",X"0004",X"0091",X"FFB6",X"FEC3",X"FEB2",X"FE41",X"FD86",X"FDA4",X"FDC9",X"FEA9",X"014F",X"03A6",X"03A1",X"02A3",X"0139",X"001C",X"FFB9",X"006B",X"007E",X"FF43",X"FEBA",X"FE91",X"FDD4",X"FD7B",X"FDA2",X"FDCD",X"FF54",X"024A",X"03A3",X"0347",X"0223",X"00CE",X"FFD3",X"FFF9",X"00BD",X"0016",X"FF18",X"FEF1",X"FE7D",X"FDC9",X"FDC0",X"FDAA",X"FE10",X"0078",X"030B",X"03A1",X"02F4",X"01A4",X"004D",X"FFAF",X"0069",X"008E",X"FF85",X"FEF3",X"FEC9",X"FDFF",X"FDA0",X"FD99",X"FD78",X"FEA0",X"01A1",X"035F",X"0394",X"028E",X"0147",X"FFE6",X"FFE5",X"00AD",X"0046",X"FF47",X"FF1A",X"FE9B",X"FDE3",X"FDC8",X"FD9C",X"FD8F",X"FFAC",X"0253",X"0387",X"0342",X"0230",X"00AB",X"FFB1",X"004C",X"00B6",X"FFB9",X"FF2A",X"FEFA",X"FE3E",X"FDCE",X"FDCF",X"FD5A",X"FE20",X"00BA",X"02D4",X"037D",X"02E3",X"01A3",X"0014",X"FFCE",X"009E",X"005D",X"FF75",X"FF46",X"FEC3",X"FE0A",X"FE05",X"FDAC",X"FD5A",X"FEFE",X"0187",X"0341",X"0370",X"02AA",X"0113",X"FFD6",X"0032",X"00BD",X"FFE8",X"FF69",X"FF1A",X"FE59",X"FDE3",X"FDF1",X"FD36",X"FDB5",X"FFE3",X"024A",X"0354",X"033F",X"0231",X"007A",X"FFDE",X"00B0",X"0083",X"FFB2",X"FF67",X"FEDB",X"FDFD",X"FE04",X"FD9A",X"FD18",X"FE46",X"00CB",X"02D9",X"0372",X"031E",X"019A",X"FFFC",X"0041",X"00D0",X"0028",X"FF9B",X"FF60",X"FE72",X"FE06",X"FE00",X"FD37",X"FD4A",X"FF12",X"019C",X"030A",X"0367",X"02A7",X"00D3",X"FFF7",X"00A9",X"009F",X"FFE3",X"FF99",X"FF1A",X"FE27",X"FE2B",X"FDBB",X"FD15",X"FDD4",X"0015",X"0241",X"0358",X"0362",X"020A",X"003C",X"003E",X"00B6",X"004A",X"FFC8",X"FF97",X"FE9A",X"FE28",X"FE19",X"FD61",X"FD11",X"FE84",X"00E9",X"02AE",X"0373",X"031E",X"012D",X"001A",X"007F",X"00AB",X"0000",X"FFF3",X"FF50",X"FE66",X"FE5A",X"FDE5",X"FD11",X"FD4F",X"FF51",X"017D",X"02E3",X"0384",X"0265",X"008D",X"0050",X"00DC",X"0086",X"0019",X"FFE9",X"FEEA",X"FE77",X"FE52",X"FD92",X"FCDD",X"FDDB",X"FFFB",X"01E3",X"0333",X"034C",X"0187",X"0033",X"0091",X"00BC",X"0033",X"002D",X"FF8D",X"FEB1",X"FE91",X"FE33",X"FD37",X"FD18",X"FE96",X"00B2",X"0264",X"0397",X"02D3",X"00EB",X"0049",X"00CB",X"007C",X"003B",X"0005",X"FF25",X"FE92",X"FE7E",X"FDC7",X"FCE8",X"FD6E",X"FF5E",X"013E",X"02FF",X"039B",X"0224",X"0079",X"00AB",X"00C0",X"005B",X"0061",X"FFAC",X"FEC3",X"FE8F",X"FE4C",X"FD5F",X"FCD4",X"FE11",X"FFFA",X"01D5",X"0379",X"0337",X"0149",X"0086",X"00DB",X"007D",X"0076",X"0030",X"FF5C",X"FEB4",X"FEAD",X"FE1F",X"FD14",X"FD2A",X"FEBA",X"006D",X"0277",X"0395",X"0270",X"00A9",X"00AE",X"009E",X"0075",X"007C",X"FFE9",X"FF03",X"FECC",X"FEA1",X"FDBC",X"FCD7",X"FDB5",X"FF3E",X"012C",X"0327",X"0380",X"01A0",X"00B3",X"00C6",X"0089",X"0086",X"005F",X"FF82",X"FEDB",X"FEC5",X"FE5F",X"FD3B",X"FD13",X"FE3F",X"FFBD",X"01EC",X"0394",X"02C6",X"010C",X"00D2",X"00A6",X"0079",X"0090",X"0024",X"FF34",X"FED4",X"FECA",X"FDF5",X"FCF4",X"FD73",X"FEA0",X"0058",X"02A7",X"038D",X"01FF",X"00F9",X"00E2",X"00A5",X"00AD",X"0099",X"FFD1",X"FF1A",X"FEFA",X"FEA6",X"FD60",X"FD00",X"FDBF",X"FF17",X"0132",X"0357",X"02F5",X"0164",X"00D8",X"00A1",X"0082",X"00AB",X"004E",X"FF74",X"FEF8",X"FF0C",X"FE38",X"FD2D",X"FD51",X"FE3B",X"FFA9",X"0233",X"0387",X"0252",X"013E",X"00E0",X"0092",X"00AD",X"00BA",X"0008",X"FF1A",X"FEFF",X"FEBE",X"FDA3",X"FD17",X"FD91",X"FE79",X"0072",X"030A",X"0327",X"01C9",X"011A",X"00C3",X"00A1",X"00D5",X"0099",X"FFAF",X"FF00",X"FF0D",X"FE53",X"FD68",X"FD37",X"FDCC",X"FEF9",X"0193",X"0353",X"0293",X"0183",X"00FB",X"00AA",X"00C4",X"00E4",X"0066",X"FF59",X"FF2F",X"FEF5",X"FDEB",X"FD31",X"FD64",X"FDE1",X"FFC5",X"0276",X"0320",X"0215",X"013F",X"00B9",X"009C",X"00D6",X"00EE",X"FFF1",X"FF3D",X"FF49",X"FEA7",X"FD94",X"FD48",X"FD7C",X"FE47",X"00E1",X"02FD",X"02C5",X"01CD",X"0102",X"009F",X"00A4",X"00F8",X"0097",X"FF98",X"FF59",X"FF2D",X"FE35",X"FD65",X"FD78",X"FD79",X"FF16",X"01DF",X"030E",X"026A",X"0192",X"00E3",X"00A0",X"00CC",X"0105",X"0024",X"FF80",X"FF63",X"FEDE",X"FDB1",X"FD6B",X"FD47",X"FDB3",X"0016",X"027F",X"02DE",X"021E",X"014A",X"00C8",X"00AE",X"010F",X"00BE",X"FFCB",X"FF73",X"FF5F",X"FE5C",X"FD83",X"FD68",X"FD35",X"FE6C",X"0136",X"02D5",X"02A0",X"01C7",X"010C",X"0095",X"00CF",X"011D",X"005F",X"FF9C",X"FF93",X"FF12",X"FDFE",X"FDAC",X"FD4A",X"FD4C",X"FF67",X"01F2",X"02C5",X"0248",X"0180",X"00C8",X"0090",X"010C",X"00ED",X"FFFF",X"FF8F",X"FF89",X"FE96",X"FDDC",X"FDAF",X"FD1A",X"FDD8",X"007E",X"0272",X"02C3",X"0217",X"0150",X"0087",X"00B9",X"011D",X"0095",X"FFB4",X"FFB4",X"FF3D",X"FE2B",X"FDC8",X"FD5C",X"FCFA",X"FEC7",X"0143",X"02A9",X"027A",X"01DF",X"00F7",X"0097",X"0116",X"012A",X"0041",X"FFD1",X"FFCC",X"FED6",X"FE0A",X"FDD6",X"FCF0",X"FD4F",X"FF9C",X"01E0",X"029C",X"0237",X"016C",X"009B",X"00AC",X"0136",X"00C2",X"FFF9",X"FFF1",X"FF78",X"FE77",X"FE2C",X"FD8F",X"FCD4",X"FE1B",X"008B",X"0251",X"0281",X"020D",X"010C",X"008F",X"00FD",X"012B",X"0057",X"FFF1",X"FFE3",X"FF05",X"FE51",X"FE1D",X"FD24",X"FD1B",X"FEF0",X"0150",X"025A",X"0263",X"01AB",X"00C2",X"00A4",X"012C",X"00DB",X"0020",X"0014",X"FFA5",X"FE9D",X"FE74",X"FDBF",X"FCDD",X"FD7A",X"FFC4",X"01B9",X"026A",X"0234",X"0145",X"0086",X"00DF",X"013E",X"0087",X"0028",X"0038",X"FF44",X"FEAC",X"FE6B",X"FD54",X"FCD0",X"FE31",X"009A",X"0204",X"0275",X"01F0",X"00E8",X"0092",X"0131",X"010A",X"0040",X"004D",X"FFE4",X"FEE3",X"FEA7",X"FE05",X"FCF9",X"FD10",X"FF28",X"013B",X"0254",X"0268",X"0199",X"0099",X"00D8",X"0134",X"008E",X"0034",X"0048",X"FF6A",X"FEE3",X"FE97",X"FDA3",X"FCB3",X"FDBB",X"FFF6",X"01AF",X"027E",X"0243",X"0110",X"008C",X"011D",X"00FE",X"0053",X"007B",X"FFFC",X"FF22",X"FEE4",X"FE69",X"FD25",X"FCD3",X"FE7E",X"0095",X"0200",X"0281",X"01CF",X"00B2",X"00D1",X"0153",X"00B0",X"0069",X"007A",X"FF9E",X"FF11",X"FEE4",X"FDE1",X"FCC3",X"FD3D",X"FF37",X"0124",X"024B",X"0270",X"0143",X"008B",X"0120",X"0116",X"007F",X"00AA",X"0033",X"FF6B",X"FF09",X"FEB9",X"FD61",X"FCB5",X"FDD7",X"FFEA",X"0196",X"0282",X"0206",X"00CF",X"00BC",X"0145",X"00BF",X"009A",X"008C",X"FFD8",X"FF31",X"FF29",X"FE56",X"FCFB",X"FD03",X"FE9E",X"0082",X"01FB",X"0272",X"0183",X"00A9",X"0121",X"0122",X"00A3",X"00C0",X"0062",X"FF88",X"FF40",X"FEFA",X"FDB6",X"FCB1",X"FD66",X"FF40",X"0101",X"0255",X"023C",X"0100",X"00CD",X"0142",X"00C7",X"00C7",X"00B8",X"000A",X"FF5F",X"FF50",X"FE9A",X"FD38",X"FCD5",X"FE13",X"FFD8",X"019A",X"0271",X"01A5",X"00B7",X"012B",X"010F",X"00C3",X"00E5",X"009D",X"FFBF",X"FF61",X"FF35",X"FE10",X"FCDC",X"FD2A",X"FEA6",X"0068",X"0216",X"0251",X"011D",X"00EF",X"0133",X"00EB",X"00CA",X"00ED",X"0041",X"FF7D",X"FF5E",X"FEDE",X"FD7A",X"FCCA",X"FDA5",X"FF4A",X"011C",X"0278",X"01E6",X"00F6",X"012C",X"010F",X"00B6",X"00D8",X"00B2",X"FFD5",X"FF70",X"FF74",X"FE7D",X"FD23",X"FD04",X"FE26",X"FFD9",X"01BF",X"0269",X"013F",X"00F4",X"0122",X"00D5",X"00CA",X"0100",X"007F",X"FFA7",X"FF9F",X"FF50",X"FDEC",X"FCF8",X"FD49",X"FE9B",X"0079",X"0235",X"01E1",X"011A",X"0126",X"010E",X"00B6",X"00F6",X"00E8",X"0021",X"FF94",X"FFA6",X"FED5",X"FD6F",X"FCF9",X"FDB3",X"FF28",X"0156",X"0240",X"0173",X"011E",X"0134",X"00DD",X"00C5",X"0119",X"0097",X"FFD6",X"FFB7",X"FF8E",X"FE4D",X"FD1A",X"FD23",X"FDFD",X"FFDB",X"01EA",X"01E9",X"012D",X"0122",X"0104",X"00B1",X"00F9",X"0103",X"0053",X"FFD0",X"FFEC",X"FF46",X"FDDA",X"FD1B",X"FD61",X"FE7B",X"00D3",X"0211",X"0185",X"0118",X"0123",X"00D6",X"00C4",X"0117",X"00D2",X"FFFD",X"FFDC",X"FFC7",X"FEB6",X"FD67",X"FD27",X"FD7F",X"FF54",X"0187",X"01EE",X"0148",X"0139",X"0117",X"00B0",X"00F5",X"0124",X"007C",X"FFE1",X"FFE5",X"FF8C",X"FE1E",X"FD3E",X"FD1B",X"FDF2",X"003B",X"01DA",X"019E",X"0124",X"0135",X"00DD",X"00BB",X"0130",X"010A",X"0039",X"FFF2",X"FFF7",X"FF1A",X"FDC3",X"FD2F",X"FD18",X"FEA5",X"00FB",X"01C2",X"0148",X"0141",X"010D",X"00BC",X"00E3",X"0158",X"00C9",X"0018",X"0014",X"FFDA",X"FE70",X"FD92",X"FD0E",X"FD75",X"FF9F",X"0179",X"0185",X"013F",X"0139",X"00E9",X"00A4",X"0135",X"013A",X"0076",X"0015",X"003E",X"FF57",X"FE19",X"FD63",X"FCF0",X"FE2B",X"0074",X"0183",X"014C",X"0139",X"010E",X"0092",X"00DA",X"014F",X"0103",X"0030",X"0035",X"000C",X"FEDD",X"FDE6",X"FD16",X"FD37",X"FF11",X"010F",X"0173",X"014E",X"0142",X"00D6",X"0093",X"011E",X"0157",X"00A5",X"0029",X"0056",X"FFA1",X"FE98",X"FD94",X"FCDE",X"FDA1",X"FFDE",X"0139",X"0148",X"0149",X"0129",X"0090",X"00B3",X"0152",X"0121",X"0058",X"0067",X"003A",X"FF4E",X"FE6A",X"FD5E",X"FCEE",X"FE82",X"0089",X"0140",X"013B",X"0150",X"00DF",X"0072",X"00DA",X"014D",X"00BB",X"004A",X"007F",X"FFD9",X"FEFF",X"FE0A",X"FCEC",X"FD5F",X"FF70",X"00F8",X"0136",X"0160",X"013A",X"00A3",X"008F",X"0140",X"013A",X"006C",X"0073",X"0044",X"FF81",X"FEB5",X"FD79",X"FCB0",X"FE05",X"000D",X"0114",X"0154",X"0178",X"010B",X"008B",X"00D6",X"0169",X"00E9",X"0069",X"0081",X"FFFE",X"FF4C",X"FE62",X"FCFC",X"FD04",X"FECD",X"0086",X"0101",X"015A",X"0157",X"00B9",X"0078",X"012E",X"014B",X"00A1",X"009B",X"0067",X"FFCD",X"FF25",X"FDDB",X"FCC0",X"FD87",X"FF98",X"00C0",X"0123",X"016F",X"0128",X"007E",X"00B0",X"0156",X"00EC",X"008B",X"00A5",X"0024",X"FFA7",X"FEBC",X"FD3F",X"FCC6",X"FE56",X"001A",X"00E5",X"015A",X"0170",X"00DA",X"005D",X"0108",X"0144",X"00AB",X"0096",X"006D",X"FFF5",X"FF79",X"FE37",X"FCD5",X"FD43",X"FF1E",X"006A",X"0119",X"0189",X"0160",X"0090",X"0097",X"012C",X"00F5",X"00A7",X"009C",X"003A",X"FFEC",X"FF31",X"FDA3",X"FCAE",X"FDE4",X"FF91",X"008A",X"012E",X"018C",X"00ED",X"0055",X"00F2",X"0143",X"00D7",X"00CE",X"0094",X"0035",X"FFE6",X"FEBF",X"FD0E",X"FCF5",X"FE94",X"FFEF",X"00BD",X"015B",X"0164",X"0084",X"007B",X"011B",X"00FF",X"00D6",X"00C9",X"006C",X"0033",X"FFB2",X"FE0D",X"FCC8",X"FD83",X"FF15",X"002C",X"00E7",X"0186",X"0106",X"0050",X"00C9",X"0122",X"00D9",X"00DF",X"009D",X"005E",X"003D",X"FF46",X"FD61",X"FCD7",X"FE11",X"FF85",X"0072",X"0152",X"0184",X"009A",X"006E",X"010B",X"00FC",X"00E3",X"00D4",X"006C",X"0052",X"001A",X"FE92",X"FCF4",X"FD3D",X"FEB4",X"FFC1",X"00A1",X"017B",X"011E",X"0064",X"00AC",X"0102",X"00F4",X"00FF",X"00A8",X"0067",X"0079",X"FFBE");
	--constant sound1 : table_type := (X"003A",X"0014",X"FFCD",X"FFB9",X"FF84",X"FFA9",X"FFAD",X"FF7F",X"FF55",X"FF5F",X"FF60",X"FF60",X"FF4C",X"FF48",X"FF3E",X"FF6B",X"FF82",X"FF92",X"FF55",X"FF32",X"FF15",X"FF14",X"FF05",X"FF36",X"FF7E",X"FF9B",X"FF98",X"FF9F",X"FFA4",X"FF8F",X"FF9B",X"FF87",X"FFA4",X"FFCB",X"FFEC",X"000F",X"0010",X"FFF9",X"FFF5",X"0009",X"0032",X"003C",X"0032",X"002C",X"0048",X"0052",X"0069",X"009B",X"00AA",X"00A0",X"00CA",X"00F0",X"0128",X"014F",X"0125",X"00ED",X"00B3",X"00A6",X"00CC",X"00EA",X"00BC",X"009E",X"0087",X"006A",X"0065",X"0018",X"0007",X"0014",X"0021",X"0016",X"FFF9",X"FFBE",X"FF6E",X"FF40",X"FF4A",X"FF50",X"FF5A",X"FF68",X"FF91",X"FF8B",X"FF66",X"FF40",X"FF5D",X"FF9F",X"FFAF",X"FF9E",X"FF7E",X"FF80",X"FF8F",X"FFB0",X"FFA1",X"FF95",X"FFF3",X"0043",X"006B",X"004D",X"0030",X"005D",X"007A",X"008E",X"0097",X"009B",X"00AB",X"00BE",X"00CE",X"00D4",X"00C4",X"00BD",X"00AC",X"009E",X"009F",X"0052",X"0017",X"0012",X"0012",X"0008",X"FFEF",X"FFD9",X"FFEF",X"FFF9",X"FFFD",X"000D",X"000A",X"FFDE",X"FFB2",X"FF8B",X"FF89",X"FF99",X"FF77",X"FF4E",X"FF4F",X"FF63",X"FF5B",X"FF31",X"FF1D",X"FF4B",X"FF4E",X"FF4A",X"FF58",X"FF6C",X"FF8E",X"FFA4",X"FF8E",X"FF85",X"FF6C",X"FF64",X"FF81",X"FF8D",X"FF8F",X"FFAA",X"FFB9",X"FFB3",X"FF94",X"FF9C",X"FFB6",X"FFE4",X"FFFC",X"001A",X"001F",X"FFFE",X"0025",X"0025",X"001D",X"003F",X"0029",X"0026",X"005A",X"006D",X"004E",X"0022",X"FFF8",X"FFE3",X"FFEB",X"FFA6",X"FF75",X"FF7E",X"FFAA",X"FFB0",X"FF7A",X"FF63",X"FF74",X"FFB0",X"FFD0",X"FFC1",X"FFA9",X"FF98",X"FFAF",X"FFE8",X"FFE4",X"FFC0",X"FF9C",X"FF9B",X"FF9E",X"FFC3",X"FFD3",X"FFEB",X"0009",X"002A",X"001C",X"0007",X"0007",X"001C",X"0013",X"FFF5",X"001A",X"0043",X"0047",X"0069",X"0072",X"0062",X"008B",X"00AF",X"00CD",X"00D8",X"00E0",X"00FC",X"011E",X"00F9",X"00E1",X"00F7",X"00C7",X"009A",X"0092",X"0072",X"0064",X"005E",X"0027",X"0001",X"FFF0",X"FFCC",X"FF71",X"FF55",X"FF64",X"FF87",X"FFB5",X"FFC4",X"FFD4",X"FFDA",X"FFBC",X"FFB0",X"FF75",X"FF65",X"FF5E",X"FF6B",X"FFB2",X"FFBA",X"FF9A",X"FF7B",X"FF4F",X"FF4A",X"FF53",X"FF89",X"FFAA",X"FFD5",X"FFED",X"0003",X"0006",X"FFE6",X"0003",X"0019",X"0059",X"007E",X"008E",X"00A8",X"00B7",X"00A3",X"009C",X"00C1",X"00D8",X"00C6",X"00C0",X"00B3",X"0095",X"0079",X"008F",X"0072",X"005F",X"005D",X"004F",X"0075",X"007A",X"005C",X"0022",X"0016",X"0022",X"0030",X"FFE0",X"FF96",X"FFD1",X"FFD9",X"FFCA",X"FFB4",X"FFE5",X"001F",X"FFF6",X"FF97",X"FF48",X"FF56",X"FF7B",X"FF92",X"FF90",X"FF7C",X"FF6C",X"FF5F",X"FF68",X"FF6B",X"FF62",X"FF78",X"FF98",X"FF88",X"FF80",X"FF79",X"FF4F",X"FF4A",X"FF57",X"FF83",X"FFAC",X"FFF4",X"002D",X"004F",X"004E",X"0018",X"0012",X"0021",X"0014",X"000D",X"0011",X"004E",X"0052",X"0037",X"0039",X"0002",X"0004",X"000F",X"FFE7",X"FFFB",X"002B",X"003C",X"FFFD",X"FFB0",X"FF7E",X"FF9F",X"FFA9",X"FF89",X"FFA3",X"FFC7",X"FFE1",X"FFEE",X"FFE6",X"FFC7",X"FFC3",X"FFEE",X"FFE0",X"FFD0",X"FFBE",X"FFD6",X"FFBB",X"FF75",X"FF33",X"FF26",X"FF34",X"FF53",X"FF4D",X"FF47",X"FF49",X"FFA9",X"000F",X"0040",X"000D",X"0020",X"0025",X"001B",X"0049",X"004E",X"005C",X"0085",X"00AC",X"00DD",X"00BF",X"00AE",X"00A6",X"0081",X"0088",X"0096",X"00AD",X"00C7",X"0093",X"0086",X"0081",X"0050",X"0066",X"0076",X"0063",X"0093",X"008F",X"0073",X"006E",X"0050",X"0011",X"FFEE",X"FFE2",X"FFE3",X"FFE4",X"FFCE",X"FFCA",X"FFB6",X"FF90",X"FF7B",X"FF7C",X"FF49",X"FF3C",X"FF6C",X"FF80",X"FFA1",X"FFC2",X"FFCA",X"FFE7",X"FFF6",X"0002",X"0002",X"0012",X"0013",X"001B",X"FFF1",X"0005",X"0013",X"003D",X"005C",X"004A",X"005E",X"0047",X"0027",X"005A",X"0087",X"007D",X"0064",X"0059",X"002F",X"0005",X"0001",X"001D",X"0029",X"0042",X"009A",X"00C0",X"00A5",X"006A",X"0006",X"FFE3",X"FFF4",X"FFFF",X"0010",X"001D",X"0016",X"0017",X"FFF3",X"FF99",X"FF88",X"FFA3",X"FF7A",X"FF7B",X"FF55",X"FF30",X"FF11",X"FEE6",X"FEF7",X"FED9",X"FEB8",X"FEDE",X"FF1E",X"FF31",X"FF27",X"FEE1",X"FEA7",X"FE91",X"FE66",X"FE6D",X"FE88",X"FEB7",X"FEDD",X"FF12",X"FF58",X"FF5C",X"FF82",X"FF86",X"FFB3",X"FFF6",X"0007",X"0023",X"0011",X"002A",X"004A",X"0077",X"0084",X"00BE",X"0104",X"010C",X"011D",X"013F",X"0138",X"011E",X"00EE",X"00D3",X"00CD",X"00F2",X"00FD",X"0103",X"0118",X"00D5",X"00E1",X"00E1",X"00A9",X"0075",X"0047",X"0042",X"0034",X"0006",X"FFF8",X"FFFB",X"FFD9",X"FFCE",X"FFD3",X"FFDA",X"FFFF",X"001A",X"0017",X"003D",X"0011",X"FFE1",X"0010",X"FFF9",X"FFC0",X"FFCE",X"FFED",X"FFF8",X"FFE9",X"FFAB",X"FF73",X"FF56",X"FF5F",X"FF7E",X"FF7A",X"FF70",X"FF71",X"FF7D",X"FF71",X"FF8A",X"FFA6",X"FFDC",X"FFF5",X"000D",X"0002",X"FFF7",X"FFF8",X"0026",X"0025",X"001E",X"0059",X"00A8",X"00BD",X"00D1",X"0106",X"0148",X"015B",X"016F",X"019C",X"0194",X"0175",X"014B",X"011F",X"00F1",X"00DD",X"00A1",X"0055",X"0000",X"FFDF",X"FFC5",X"FF76",X"FF45",X"FF0D",X"FEFB",X"FED7",X"FE97",X"FE3A",X"FDFF",X"FDFE",X"FE04",X"FE0C",X"FDDE",X"FDDE",X"FDFE",X"FE45",X"FE87",X"FE6B",X"FEE3",X"FF67",X"0024",X"00B5",X"010C",X"018B",X"01CD",X"0204",X"01EB",X"01EE",X"0207",X"01EB",X"01CB",X"0185",X"00FC",X"0094",X"0054",X"FFF6",X"FF8D",X"FF5A",X"FF46",X"FF35",X"FEE5",X"FE62",X"FE42",X"FE09",X"FDC6",X"FD66",X"FCF8",X"FCB5",X"FCC5",X"FCBC",X"FCB8",X"FD28",X"FDEC",X"FECE",X"FFD2",X"00E9",X"024B",X"0395",X"04A2",X"051D",X"055B",X"05A9",X"0584",X"04F2",X"03FC",X"02F2",X"0208",X"0118",X"FFE9",X"FEC0",X"FDCD",X"FD10",X"FC7F",X"FC23",X"FBC7",X"FBA7",X"FB89",X"FB77",X"FB78",X"FB5C",X"FAF3",X"FB02",X"FAC4",X"FAF1",X"FBB8",X"FC9B",X"FE04",X"FF51",X"0153",X"035F",X"054E",X"075B",X"08DD",X"09D2",X"0A1B",X"0995",X"0877",X"0718",X"0612",X"0420",X"02C1",X"017E",X"FFF2",X"FF26",X"FE03",X"FD2A",X"FC4E",X"FC14",X"FC2E",X"FC29",X"FC5B",X"FC85",X"FCFD",X"FD07",X"FC98",X"FC0E",X"FB0D",X"FA6C",X"F98F",X"F97B",X"F9EF",X"FAA3",X"FC9B",X"FE50",X"011A",X"0386",X"05FE",X"0837",X"0972",X"0A3A",X"0A64",X"0931",X"0788",X"051C",X"03EC",X"0295",X"0149",X"002E",X"FEEC",X"FEB0",X"FE64",X"FDD2",X"FD60",X"FD05",X"FD0E",X"FD5F",X"FD39",X"FD1D",X"FD53",X"FD4E",X"FC93",X"FB40",X"FA02",X"F8D9",X"F808",X"F895",X"F913",X"F9F8",X"FBEA",X"FE76",X"0261",X"057B",X"094A",X"0AE3",X"0C84",X"0CFA",X"0C82",X"0ABD",X"072E",X"03CC",X"004B",X"FDF6",X"FDCB",X"FD0C",X"FC89",X"FDA6",X"FE89",X"FFBC",X"FF7C",X"FF1A",X"FF39",X"FF68",X"FF21",X"FDFD",X"FD1F",X"FC5C",X"FB6B",X"F9AF",X"F79F",X"F5D5",X"F4C4",X"F405",X"F52A",X"F5F9",X"F7C4",X"FA75",X"FE6A",X"0330",X"085B",X"0BD0",X"0E21",X"0FD0",X"1035",X"0FF4",X"0C69",X"0811",X"0343",X"003B",X"FEA8",X"FCDD",X"FCB0",X"FC60",X"FDF9",X"FF18",X"FF55",X"FFA8",X"FFB1",X"00BC",X"00C6",X"002C",X"FF37",X"FE5D",X"FD8E",X"FBD6",X"F965",X"F6CB",X"F505",X"F3AC",X"F366",X"F486",X"F5B6",X"F824",X"FB81",X"008E",X"0730",X"0C3A",X"0EEA",X"1135",X"11C5",X"1243",X"0F5E",X"0A82",X"04DE",X"00AA",X"FE9E",X"FC69",X"FA5D",X"F9AE",X"FA92",X"FCBF",X"FDD6",X"FE1D",X"FEBB",X"FFED",X"013A",X"012E",X"0014",X"FF52",X"FE98",X"FD06",X"FA86",X"F786",X"F530",X"F388",X"F24C",X"F308",X"F44E",X"F69B",X"F9DB",X"FF3B",X"066F",X"0C2A",X"100F",X"131D",X"1413",X"154C",X"12ED",X"0E90",X"08A9",X"03C8",X"0123",X"FE16",X"FB8E",X"F9D2",X"FA0A",X"FB9C",X"FC52",X"FC81",X"FCF9",X"FE7A",X"FFBB",X"FFB0",X"FF44",X"FE82",X"FD59",X"FBCD",X"F924",X"F620",X"F444",X"F19D",X"EFAB",X"EFD1",X"F1C5",X"F49B",X"F886",X"FD96",X"0495",X"0C54",X"10B0",X"14B6",X"155B",X"1625",X"149D",X"0FF1",X"09C8",X"0367",X"FF17",X"FC28",X"FB3B",X"F9CD",X"F9E1",X"FC02",X"FD29",X"FF76",X"FF2B",X"FF56",X"FFAC",X"002A",X"00AE",X"FF0E",X"FD92",X"FB82",X"F9A5",X"F7CA",X"F449",X"F107",X"EE9D",X"EE9C",X"F062",X"F1FC",X"F514",X"FAA6",X"0498",X"0C10",X"1200",X"154F",X"164F",X"186A",X"1699",X"12B0",X"0B33",X"04C4",X"00E4",X"FDB0",X"FAD6",X"F7F8",X"F6F9",X"F923",X"FB64",X"FC9B",X"FCAA",X"FDA0",X"FF17",X"0030",X"FFCB",X"FED6",X"FE92",X"FD1B",X"FAB1",X"F71F",X"F471",X"F0B3",X"EE00",X"EE80",X"F04A",X"F2F6",X"F6F6",X"FDEB",X"08B0",X"0EA1",X"1477",X"17F6",X"197E",X"1A6C",X"181E",X"1171",X"09CB",X"031F",X"FF3A",X"FBDB",X"F8DD",X"F746",X"F874",X"FB03",X"FCF9",X"FD8C",X"FE62",X"FF50",X"FFB4",X"004F",X"FF54",X"FDE3",X"FCD9",X"FA5B",X"F7A9",X"F378",X"F109",X"EDDB",X"EBEF",X"ED80",X"F051",X"F4BD",X"FBF5",X"0718",X"1034",X"166D",X"195F",X"1897",X"19C1",X"1678",X"10BD",X"0903",X"0130",X"FD7C",X"FAC4",X"F8A8",X"F7A3",X"F894",X"FC0B",X"FFD3",X"00F3",X"01A1",X"0359",X"02EE",X"022C",X"0069",X"FDC0",X"FCB5",X"FA29",X"F6EF",X"F371",X"EFEF",X"EE0B",X"ECF4",X"EE12",X"F397",X"F8AF",X"FE30",X"08B4",X"1392",X"16E1",X"19CB",X"15F4",X"1294",X"1111",X"08E3",X"FF7D",X"F883",X"F692",X"FAA3",X"FC66",X"FE81",X"0361",X"072A",X"09AD",X"0753",X"0107",X"FDA4",X"FBC1",X"F885",X"F7BF",X"F713",X"F8F3",X"F9E9",X"F778",X"F5B9",X"F007",X"EEB3",X"EAA0",X"EB52",X"F525",X"F8A0",X"0305",X"10EB",X"1C75",X"2156",X"1F40",X"1383",X"09FF",X"01E9",X"F76F",X"EF4B",X"EA84",X"F257",X"0309",X"0B5B",X"1446",X"169E",X"145E",X"10B1",X"0245",X"F494",X"EF3F",X"ECEF",X"F1B1",X"F7B8",X"FB20",X"00DE",X"0231",X"FDF6",X"F977",X"EE32",X"E9E1",X"E4E8",X"E02D",X"EE2E",X"F7D0",X"04C9",X"19CE",X"2799",X"27D3",X"2217",X"0E31",X"FECD",X"F5DA",X"EB6E",X"E820",X"EC8D",X"FCA4",X"1216",X"1AEB",X"1E35",X"187A",X"0D07",X"024C",X"F23C",X"E96D",X"ECED",X"F489",X"FF2B",X"058B",X"06D2",X"0706",X"01DD",X"F841",X"F1D2",X"E9DC",X"E839",X"E5EA",X"E7CA",X"F7EB",X"0599",X"13CA",X"27AB",X"2609",X"1CD8",X"10E6",X"FB89",X"EF9E",X"EB78",X"E588",X"F02D",X"FED6",X"13EA",X"2245",X"2227",X"18D4",X"0ACC",X"F9FE",X"ED9F",X"E559",X"E97B",X"F79B",X"0374",X"09F5",X"09FF",X"0639",X"0045",X"F7D1",X"EF15",X"EB21",X"E83C",X"E6A4",X"E5F5",X"F2BD",X"03F2",X"1377",X"228C",X"2799",X"1C01",X"10A2",X"FE2B",X"ED8D",X"E996",X"E861",X"F0E2",X"0019",X"159A",X"23B1",X"2369",X"179A",X"074E",X"F6DD",X"ECCA",X"E696",X"EC13",X"FA38",X"06FF",X"0B94",X"095F",X"0360",X"FD4E",X"F5FC",X"EE4B",X"EB05",X"EB23",X"EB55",X"E69C",X"F03A",X"0414",X"1162",X"1D9A",X"26E2",X"1B84",X"0FD8",X"FE50",X"ED07",X"E907",X"EA76",X"F0C0",X"006D",X"14AE",X"23BD",X"2342",X"1650",X"0516",X"F422",X"EBD6",X"E823",X"EE45",X"FCA0",X"0924",X"0D2C",X"0874",X"018D",X"FC15",X"F49E",X"EF52",X"EC7B",X"EB6A",X"ED6C",X"E9FD",X"EF1D",X"023B",X"0D53",X"1958",X"285D",X"1E0A",X"0FDA",X"00E2",X"EF18",X"E9A9",X"EC2F",X"EFC5",X"FF47",X"1514",X"2326",X"22B4",X"1542",X"038C",X"F416",X"EC34",X"E949",X"EFDA",X"FCE4",X"0903",X"0C72",X"071D",X"FFCE",X"FA35",X"F530",X"F002",X"EEB7",X"ED76",X"EB1A",X"E6AB",X"ECCA",X"028B",X"11D7",X"1E33",X"2B26",X"2004",X"10C1",X"FFE6",X"ECA8",X"E755",X"EB09",X"F234",X"0437",X"1999",X"265C",X"248F",X"1470",X"007C",X"EFBA",X"E8ED",X"E8C2",X"F2DB",X"00CD",X"0C79",X"0EBE",X"0710",X"FEC2",X"F8B1",X"F3C8",X"EFA8",X"ED6E",X"EBEE",X"EBDB",X"E70B",X"EF88",X"046C",X"13FB",X"2347",X"2AE4",X"1B90",X"0CF8",X"FA67",X"E92B",X"E6DB",X"EA35",X"F4E7",X"08D7",X"1D3C",X"27A3",X"2204",X"0E2E",X"FA2B",X"EAAF",X"E64E",X"EA85",X"F67D",X"0455",X"0EE3",X"0EFD",X"050D",X"FBE6",X"F502",X"F131",X"EDC4",X"EE4C",X"ECE3",X"E99E",X"E434",X"F2B6",X"094C",X"1A04",X"2A0E",X"2928",X"15B2",X"080A",X"F4C4",X"E627",X"E773",X"EC32",X"FB0D",X"10B7",X"232A",X"28C1",X"1EB0",X"089C",X"F361",X"E71D",X"E5DD",X"EDFB",X"FB57",X"08E6",X"0F8D",X"0C73",X"003D",X"F92C",X"F436",X"F165",X"EDFC",X"EBF0",X"EA12",X"E6FE",X"E59A",X"F8FC",X"0E4C",X"1F30",X"2E07",X"249C",X"0F9F",X"FF82",X"ED03",X"E38B",X"E791",X"EFA6",X"023A",X"197D",X"289C",X"2789",X"1859",X"FFC3",X"ECC2",X"E6E1",X"E7F9",X"F39B",X"01CF",X"0BED",X"0F47",X"08AA",X"FCE4",X"F861",X"F50F",X"F314",X"F1BF",X"EE0C",X"EA4F",X"E419",X"E833",X"FE54",X"12CE",X"22E5",X"2E43",X"1F10",X"0CBA",X"F9EA",X"E80E",X"E50B",X"EA75",X"F418",X"089D",X"1EDE",X"29E4",X"251E",X"10A7",X"F84C",X"E94C",X"E5C0",X"EB35",X"F90C",X"055F",X"0DB4",X"0D6A",X"02E2",X"FA8A",X"F715",X"F4B0",X"F336",X"F09A",X"EC80",X"E8A9",X"E1E4",X"EF52",X"0641",X"18DF",X"29F7",X"2AE0",X"15FE",X"05D1",X"F1C7",X"E419",X"E70E",X"EE3F",X"FC0E",X"1312",X"2585",X"298F",X"1FB0",X"0776",X"F15F",X"E886",X"E8B9",X"F319",X"018F",X"0A4B",X"0EF4",X"0B47",X"FEB6",X"F94B",X"F655",X"F44F",X"F316",X"EFA1",X"ED23",X"E914",X"E4B3",X"F5D2",X"0B07",X"1BDB",X"2D28",X"25F5",X"0EE6",X"FDC9",X"EBE4",X"E388",X"E88D",X"EFB7",X"FFE1",X"1780",X"26E4",X"26C4",X"1848",X"FEC5",X"EBFF",X"E6B2",X"EA83",X"F777",X"0382",X"0AFB",X"0CD3",X"0505",X"FA83",X"F60C",X"F3DD",X"F3BF",X"F313",X"F02F",X"ECD3",X"E625",X"E838",X"FB39",X"0FE6",X"21B6",X"2DC7",X"20A7",X"0C99",X"F905",X"E88F",X"E499",X"EA32",X"F46F",X"08F0",X"1F20",X"295A",X"246D",X"0FAB",X"F722",X"E980",X"E869",X"F09D",X"FEAC",X"088C",X"0D6F",X"0B5D",X"0138",X"F8F6",X"F5A0",X"F4CB",X"F4EB",X"F39F",X"EEDE",X"EA12",X"E394",X"EDE8",X"032D",X"1720",X"2660",X"294B",X"177D",X"061E",X"F1BD",X"E400",X"E500",X"EC45",X"F903",X"1020",X"227C",X"270C",X"1DE9",X"0645",X"F0C0",X"E85C",X"E999",X"F4BC",X"019E",X"08F1",X"0BA6",X"0692",X"FCA6",X"F894",X"F691",X"F71C",X"F614",X"F30B",X"EDE8",X"E80D",X"E4A4",X"F4A2",X"09DF",X"1E08",X"2D85",X"2944",X"1400",X"00C1",X"ED4C",X"E3FD",X"E776",X"EFE7",X"FFDE",X"16FF",X"26F2",X"2799",X"17EB",X"0010",X"ED7F",X"E7E1",X"ED74",X"FA6E",X"046D",X"0A86",X"09E7",X"024D",X"FAAB",X"F854",X"F72B",X"F767",X"F476",X"EFBF",X"E9B6",X"E4B2",X"E8EE",X"FB72",X"0F92",X"2227",X"2C9B",X"2090",X"0CE7",X"F74F",X"E68D",X"E40D",X"E9E0",X"F4BD",X"08F5",X"1CC3",X"2563",X"2121",X"0DB1",X"F76A",X"EB6C",X"EA5E",X"F290",X"FEC4",X"0634",X"0975",X"0759",X"0054",X"FBA7",X"FA07",X"F885",X"F694",X"F348",X"ED45",X"E815",X"E405",X"F184",X"05CF",X"1995",X"2A4C",X"2A77",X"1758",X"0561",X"F022",X"E47C",X"E6B3",X"EE06",X"FBB0",X"1194",X"2210",X"258F",X"1B05",X"046D",X"F081",X"E8F8",X"EBFD",X"F6D3",X"014E",X"076D",X"0830",X"03B5",X"FC81",X"F9F2",X"F838",X"F69F",X"F465",X"F0C2",X"E9C3",X"E4FF",X"E649",X"F68B",X"0A49",X"1D83",X"2C16",X"24B0",X"10BE",X"FCE5",X"EB05",X"E564",X"EA1A",X"F308",X"03BC",X"1734",X"23D2",X"22FF",X"12C1",X"FCF5",X"ED98",X"E999",X"F0E1",X"FCF0",X"0537",X"0990",X"07D2",X"0143",X"FBAB",X"F9D5",X"F97F",X"F770",X"F4A9",X"F052",X"EA1E",X"E56A",X"EF26",X"FFB0",X"1109",X"2158",X"2977",X"1D3B",X"0B5B",X"F5EF",X"E7E8",X"E769",X"EE23",X"F83F",X"0A1C",X"1A45",X"222C",X"1D1D",X"0AB0",X"F63A",X"EBC8",X"EC4F",X"F537",X"FFEA",X"066F",X"07F2",X"04E6",X"FDD3",X"FA94",X"F9A7",X"F867",X"F590",X"F2F2",X"EC8D",X"E85D",X"E63D",X"F269",X"049D",X"17D2",X"25FC",X"2725",X"166D",X"0572",X"F1FA",X"E77A",X"E982",X"F1BE",X"FDF6",X"117D",X"1FE1",X"2329",X"1904",X"04AA",X"F20B",X"EBCD",X"EFDA",X"FAAB",X"0434",X"090C",X"08CF",X"03FD",X"FCFB",X"FAB0",X"F9B9",X"F91E",X"F710",X"F387",X"ECAF",X"E8EF",X"E8EA",X"F5FF",X"06DD",X"1940",X"278B",X"23F8",X"1212",X"0061",X"EDF6",X"E6E6",X"EAFE",X"F355",X"01F3",X"144A",X"1F34",X"1FBA",X"11E7",X"FC97",X"ED9E",X"E969",X"EFDB",X"FC2E",X"0403",X"07C3",X"05CF",X"FF71",X"FAB3",X"F949",X"F86E",X"F762",X"F4FA",X"F041",X"E981",X"E591",X"EC97",X"FCCC",X"0CD7",X"1D15",X"278B",X"209E",X"0EED",X"FC0D",X"EC39",X"E85B",X"EE6F",X"F891",X"09C2",X"1ACE",X"217A",X"1DA9",X"0D36",X"F8FF",X"EE91",X"EDC9",X"F554",X"FF9A",X"055C",X"06E8",X"03D3",X"FDB7",X"FAF9",X"F950",X"F7AA",X"F639",X"F3CA",X"EF74",X"EB28",X"E68B",X"EE7F",X"FEF7",X"0EF7",X"1D6D",X"25C2",X"1B6A",X"0A20",X"F78E",X"EA7D",X"E8EF",X"EF20",X"F85E",X"0A2A",X"1962",X"1F19",X"1A48",X"08B6",X"F6C1",X"EE5B",X"EE3A",X"F6C0",X"FFF1",X"04EF",X"06E5",X"0339",X"FD0F",X"FAC3",X"F9A8",X"F948",X"F6F2",X"F439",X"EFAD",X"EC10",X"E9EB",X"F381",X"02AB",X"1362",X"1F61",X"2562",X"1AA0",X"0900",X"F5C0",X"EA8B",X"EA68",X"F24F",X"FCBB",X"0EE3",X"1C0D",X"2138",X"1916",X"05B6",X"F4FE",X"EEB8",X"F09F",X"F9D4",X"01C8",X"064E",X"0671",X"026E",X"FCFA",X"FA78",X"F857",X"F7F6",X"F5A4",X"F336",X"EEA5",X"EB00",X"E912",X"F3FB",X"03F4",X"143D",X"1F5D",X"21BD",X"153F",X"0602",X"F3C2",X"EA58",X"EB83",X"F2FD",X"FEB3",X"1105",X"1C54",X"1E57",X"1461",X"0267",X"F415",X"EF15",X"F1AA",X"FB4B",X"026C",X"0618",X"060B",X"017A",X"FC9E",X"FAE9",X"F941",X"F921",X"F6BB",X"F400",X"F036",X"EBE4",X"EA51",X"F563",X"04AB",X"14EE",X"1FAC",X"2104",X"15CC",X"0588",X"F3E1",X"EB57",X"EC5C",X"F388",X"FF7E",X"10B0",X"1C67",X"1E7C",X"1447",X"01A1",X"F2AD",X"ED92",X"F07E",X"F9CC",X"0180",X"0591",X"05DF",X"0147",X"FBFC",X"FA05",X"F83A",X"F78C",X"F499",X"F151",X"ECD8",X"E833",X"E7E5",X"F421",X"0485",X"1517",X"2036",X"2195",X"1677",X"05BC",X"F305",X"E96D",X"EAEB",X"F339",X"00A3",X"12F3",X"1DC0",X"1E9C",X"13DA",X"004D",X"F28C",X"EE6B",X"F19F",X"FB1A",X"01B1",X"0568",X"0590",X"0116",X"FD40",X"FB88",X"F9B3",X"F8C6",X"F5D4",X"F26D",X"EE04",X"E8AB",X"E938",X"F62C",X"0711",X"161D",X"1FBA",X"2104",X"1656",X"05A9",X"F3C3",X"EA51",X"EBF9",X"F423",X"01B1",X"139E",X"1DE7",X"1E68",X"12CE",X"0032",X"F3ED",X"EFAF",X"F2E0",X"FC20",X"021A",X"05C7",X"0655",X"01A0",X"FD9F",X"FBA4",X"F9F7",X"F934",X"F601",X"F221",X"ED65",X"E883",X"E969",X"F67C",X"07B4",X"1633",X"1F18",X"202C",X"158D",X"05A5",X"F4DE",X"EB0D",X"EC64",X"F4FC",X"02A9",X"14BF",X"1EE6",X"1E98",X"130F",X"0054",X"F3C1",X"F00D",X"F2C0",X"FBD9",X"021F",X"05B4",X"0687",X"0255",X"FDD4",X"FB77",X"F8D3",X"F77D",X"F413",X"F0DE",X"EDEB",X"EA76",X"EB5A",X"F6C8",X"064D",X"1421",X"1B8D",X"1CD5",X"144D",X"0479",X"F49D",X"EC44",X"ED12",X"F58A",X"0323",X"13E3",X"1CAE",X"1C55",X"0FD4",X"FDBD",X"F352",X"F03C",X"F363",X"FCD4",X"02DD",X"0603",X"0615",X"0139",X"FCAF",X"F9C9",X"F812",X"F750",X"F401",X"F17E",X"EE4C",X"EA54",X"EB66",X"F71B",X"05B9",X"12C1",X"1B26",X"1BCD",X"12C7",X"04D6",X"F585",X"ED73",X"EF25",X"F6C7",X"03A6",X"132C",X"1B5F",X"1B3D",X"0E95",X"FD6C",X"F36B",X"F03A",X"F490",X"FDF3",X"038A",X"06F1",X"0633",X"0007",X"FA3C",X"F738",X"F65D",X"F6C9",X"F497",X"F17D",X"ECB6",X"E90E",X"EC9C",X"F96A",X"07C3",X"14BE",X"1C5D",X"1C30",X"137B",X"04CD",X"F452",X"EC08",X"EE05",X"F70C",X"05DD",X"163C",X"1C6A",X"1ABE",X"0D4D",X"FB6F",X"F210",X"F02E",X"F590",X"FEC3",X"03E7",X"0743",X"05AF",X"FFA1",X"FB14",X"F819",X"F74F",X"F795",X"F47A",X"F1FD",X"EDF8",X"E9E3",X"EDB5",X"F90E",X"071A",X"154F",X"1CAE",X"1D18",X"1511",X"05A0",X"F675",X"EE77",X"EF65",X"F832",X"068B",X"165B",X"1DC9",X"1B5F",X"0DCC",X"FCC5",X"F2FE",X"F1B2",X"F6BE",X"FF04",X"03E6",X"0634",X"049B",X"FF3B",X"FA9D",X"F7BD",X"F76F",X"F7C1",X"F5C9",X"F29F",X"ED9D",X"E955",X"EE51",X"FA04",X"07BE",X"1437",X"1C37",X"1C94",X"1496",X"04E5",X"F51C",X"EC77",X"EE44",X"F708",X"06B2",X"1640",X"1C98",X"1AD6",X"0D19",X"FB62",X"F247",X"F056",X"F5EA",X"FE43",X"02CB",X"05ED",X"0452",X"FECD",X"FA9A",X"F779",X"F731",X"F662",X"F486",X"F2D7",X"EDD2",X"E948",X"EDA4",X"F95D",X"06DF",X"1350",X"1CC1",X"1CF1",X"13B8",X"04A9",X"F4A7",X"EC60",X"EF06",X"F721",X"06F8",X"1689",X"1BD9",X"198C",X"0BDB",X"FAEE",X"F2C1",X"F16E",X"F740",X"FEE3",X"02DD",X"04FE",X"02A5",X"FD87",X"FA0C",X"F762",X"F753",X"F6F6",X"F420",X"F19D",X"ED3E",X"E9D0",X"F002",X"FC2E",X"08D4",X"1528",X"1CF7",X"1BDF",X"1294",X"02C0",X"F3D7",X"ED3C",X"F047",X"F968",X"093B",X"183D",X"1D1B",X"1843",X"0A01",X"F93E",X"F07B",X"F0EA",X"F7C2",X"FF8D",X"0436",X"05AC",X"0344",X"FDDA",X"F960",X"F757",X"F765",X"F633",X"F407",X"F0BA",X"ED00",X"EB39",X"F0F6",X"FCCF",X"08FF",X"1480",X"1CD8",X"1B7F",X"122A",X"0308",X"F44F",X"EE53",X"F1D0",X"FAE1",X"0B6F",X"187E",X"1BD7",X"1702",X"08E7",X"FA5C",X"F305",X"F2E6",X"F9B3",X"FFA6",X"0318",X"04A8",X"0222",X"FE00",X"FAD8",X"F8F2",X"F8C2",X"F67B",X"F3B5",X"F0C1",X"ECC3",X"EB72",X"F157",X"FD9C",X"0A3C",X"1520",X"1C5A",X"1A7D",X"10FE",X"0228",X"F47F",X"EF0F",X"F236",X"FB12",X"0B54",X"1962",X"1CEF",X"1658",X"0785",X"F8EA",X"F196",X"F1F5",X"F8AA",X"FF03",X"02D7",X"03C1",X"011A",X"FCD9",X"F98F",X"F81F",X"F845",X"F6DB",X"F482",X"F091",X"ED07",X"EB2F",X"F07C",X"FD59",X"0A9E",X"15D2",X"1DBD",X"1AF4",X"104E",X"00F2",X"F2F0",X"EE3E",X"F26D",X"FC64",X"0D89",X"197E",X"1BB5",X"14B1",X"055D",X"F86E",X"F2C4",X"F374",X"FA97",X"0000",X"0315",X"0391",X"0016",X"FBFF",X"F9A3",X"F8A8",X"F871",X"F5D8",X"F309",X"EF11",X"EBBF",X"EA70",X"F0EC",X"FE45",X"0B99",X"1653",X"1CCE",X"195E",X"0E21",X"FEC0",X"F1D9",X"EDD7",X"F2C7",X"FD60",X"0E11",X"1946",X"1B3F",X"1315",X"038D",X"F7C4",X"F2F5",X"F3D9",X"FAC3",X"FF90",X"0271",X"02D5",X"FF47",X"FB8F",X"F96E",X"F87D",X"F83B",X"F639",X"F359",X"EF53",X"EBB5",X"EA9A",X"F3AF",X"01F4",X"0DF9",X"185F",X"1D18",X"176F",X"0BD4",X"FCEF",X"F1CC",X"EFC0",X"F51D",X"0110",X"1097",X"1993",X"1A21",X"1089",X"015B",X"F70C",X"F3CE",X"F69E",X"FCD4",X"00D9",X"02BA",X"01B0",X"FF00",X"FC08",X"FA86",X"FA36",X"F87F",X"F590",X"F233",X"ED99",X"EB7F",X"EC9A",X"F65C",X"055D",X"1190",X"19F1",X"1BF4",X"146A",X"0776",X"F9A1",X"F114",X"F144",X"F786",X"05A5",X"141E",X"199F",X"188B",X"0D74",X"FE6B",X"F68B",X"F46E",X"F8BC",X"FE6B",X"00FA",X"02C9",X"0163",X"FDBA",X"FAE8",X"F975",X"F9D0",X"F8E7",X"F545",X"F11F",X"EDD8",X"EBC2",X"EEFE",X"FADC",X"07C6",X"129E",X"1AE1",X"1A6D",X"11C7",X"03BC",X"F5D4",X"EF5D",X"F14B",X"F936",X"093E",X"16AE",X"1A76",X"14B7",X"07D0",X"FAFA",X"F4CB",X"F573",X"FB19",X"FFC1",X"0233",X"0298",X"004A",X"FD18",X"FA99",X"F9AA",X"F8CF",X"F784",X"F544",X"F0AD",X"ED01",X"EB80",X"F204",X"FF11",X"0BEB",X"15EC",X"1BAB",X"1759",X"0C91",X"FE13",X"F247",X"EEE3",X"F347",X"FEE9",X"0EEF",X"1836",X"19A3",X"101F",X"010E",X"F79E",X"F39E",X"F622",X"FCC6",X"0092",X"02DC",X"0231",X"FECD",X"FBED",X"FA5C",X"FA00",X"F8BD",X"F645",X"F3C8",X"EFE0",X"EC87",X"ED72",X"F6E9",X"0467",X"1025",X"189F",X"1A76",X"13B1",X"06F9",X"F924",X"F03E",X"EF99",X"F604",X"052B",X"1373",X"18F8",X"1640",X"0A67",X"FB9A",X"F467",X"F3FB",X"F8CD",X"FE81",X"0172",X"023E",X"00C0",X"FDB7",X"FAD9",X"FA1D",X"F9C4",X"F741",X"F4B3",X"F160",X"EE75",X"EBDA",X"F013",X"FC47",X"0994",X"1451",X"1B8E",X"193A",X"0FE9",X"0186",X"F536",X"F022",X"F359",X"FCD6",X"0C9A",X"17C6",X"19BA",X"1219",X"0437",X"F990",X"F5C5",X"F710",X"FC8F",X"0037",X"0156",X"005F",X"FDEC",X"FB28",X"FA75",X"FB21",X"FB1D",X"F7BD",X"F39E",X"EF16",X"EB7A",X"EBDD",X"F48F",X"023C",X"0F66",X"18B7",X"1C34",X"16D0",X"0ACA",X"FC6B",X"F260",X"F071",X"F5D4",X"033E",X"1218",X"18D2",X"17CD",X"0D58",X"FEF6",X"F714",X"F56C",X"F90B",X"FE33",X"00D3",X"0168",X"FFDC",X"FCDD",X"FB03",X"FB32",X"FC17",X"FA22",X"F60C",X"F18A",X"ED59",X"EB15",X"EEBA",X"FA33",X"074A",X"126D",X"1AFB",X"1AC7",X"126F",X"046F",X"F641",X"EFCF",X"F27B",X"FAE5",X"0AD9",X"16FA",X"1975",X"1296",X"0568",X"FA70",X"F5C5",X"F673",X"FBE5",X"FF54",X"008D",X"0022",X"FD1F",X"FA76",X"F9FF",X"FA94",X"FA54",X"F77D",X"F3DE",X"EF28",X"EB14",X"EABF",X"F2FA",X"00BD",X"0E2A",X"17EE",X"1BDC",X"16C2",X"0AFD",X"FC5D",X"F201",X"F00C",X"F566",X"028D",X"1168",X"182A",X"179E",X"0DAD",X"FEF4",X"F71A",X"F629",X"F97F",X"FE4B",X"FFE9",X"FFD8",X"FE5A",X"FBD4",X"FAAA",X"FAF7",X"FB86",X"F96D",X"F51F",X"F0C7",X"EBBE",X"E928",X"EE16",X"F9C4",X"0746",X"128A",X"1AEB",X"1AD4",X"120D",X"0402",X"F67C",X"EFF5",X"F20D",X"FA97",X"0AA7",X"16E2",X"1960",X"12AF",X"05EF",X"FB6D",X"F707",X"F7B7",X"FD02",X"0040",X"00C3",X"0058",X"FDAF",X"FBAE",X"FBB3",X"FC6B",X"FC5B",X"F8B0",X"F429",X"EE8B",X"EB45",X"EB8B",X"F335",X"00A4",X"0D57",X"16C7",X"1BD9",X"174C",X"0BDC",X"FD29",X"F280",X"F075",X"F5FD",X"039E",X"1257",X"1769",X"1590",X"0C10",X"FF45",X"F8B5",X"F7D6",X"FACD",X"FEAC",X"FFF8",X"FFB5",X"FDF9",X"FBEF",X"FB0F",X"FB9D",X"FD1F",X"FB59",X"F694",X"F283",X"EDD4",X"EB02",X"EF0F",X"F9B5",X"0696",X"1216",X"19F1",X"19B1",X"11BB",X"03B7",X"F70E",X"F137",X"F31A",X"FB5A",X"0A58",X"1567",X"17F1",X"108B",X"044E",X"FB98",X"F7F7",X"F98D",X"FEC4",X"0111",X"00D8",X"FF18",X"FBE0",X"FA67",X"FB17",X"FCD2",X"FD1F",X"F951",X"F502",X"EFEF",X"EC38",X"EBF7",X"F39D",X"001D",X"0CD4",X"158D",X"19EA",X"15C2",X"0AD5",X"FCC4",X"F346",X"F197",X"F71A",X"0435",X"1124",X"1516",X"128A",X"096A",X"FE24",X"F87E",X"F7E4",X"FB94",X"FF48",X"FF9F",X"FECB",X"FCD3",X"FB01",X"FA5C",X"FB4A",X"FC96",X"FB02",X"F6AC",X"F259",X"ED81",X"EB66",X"F03E",X"FAB1",X"05D9",X"0FFE",X"16D9",X"1755",X"104E",X"0371",X"F7B3",X"F287",X"F40E",X"FC5D",X"0B10",X"13F4",X"154A",X"0D56",X"0174",X"FA9F",X"F805",X"F98F",X"FE9A",X"0014",X"0038",X"FECC",X"FBC4",X"FAB0",X"FB0E",X"FC87",X"FCBC",X"F91F",X"F4F0",X"F126",X"ED91",X"ECD3",X"F462",X"00ED",X"0D08",X"1525",X"18EF",X"14B3",X"0A89",X"FD76",X"F4D5",X"F344",X"F84C",X"054F",X"1187",X"1436",X"10E6",X"06E0",X"FCB1",X"F8AD",X"F8BF",X"FCEE",X"00AD",X"00CF",X"FF8F",X"FCE6",X"FA9F",X"FA80",X"FC27",X"FDC7",X"FB94",X"F727",X"F398",X"EEF1",X"ECD3",X"F231",X"FC0B",X"06C0",X"1190",X"1861",X"17A0",X"1014",X"03F0",X"F964",X"F465",X"F5F3",X"FE07",X"0C2F",X"14BE",X"1513",X"0D45",X"01D0",X"FB04",X"F970",X"FB10",X"0009",X"015B",X"008C",X"FEFE",X"FBCB",X"FA5A",X"FB18",X"FC6D",X"FC5F",X"F92F",X"F4ED",X"F029",X"ECE2",X"EC5A",X"F3EC",X"00AD",X"0BF7",X"1423",X"1878",X"1486",X"0B60",X"FEE8",X"F5EE",X"F3AF",X"F7A2",X"02D6",X"0FD1",X"13DD",X"1255",X"08DF",X"FD6F",X"F976",X"F965",X"FBEE",X"FF42",X"FF10",X"FE5F",X"FC74",X"FA37",X"FA54",X"FBB5",X"FCBA",X"FB00",X"F615",X"F22B",X"EEA8",X"EC0C",X"EE6C",X"F7C9",X"03A2",X"0E9D",X"164A",X"1763",X"1149",X"06AE",X"FB92",X"F520",X"F565",X"FA7F",X"0788",X"1293",X"1439",X"0F20",X"0521",X"FC1C",X"F991",X"FA31",X"FE10",X"FFF5",X"FEE0",X"FE0D",X"FC5A",X"FB19",X"FBFD",X"FD1C",X"FD41",X"FA04",X"F50A",X"F108",X"EEAF",X"ED87",X"F118",X"FAE3",X"063E",X"109C",X"180C",X"16EC",X"0FA3",X"03E9",X"F9DA",X"F59D",X"F741",X"FE2F",X"0B4E",X"1345",X"1430",X"0CE9",X"023F",X"FC45",X"FAD2",X"FBDB",X"FF36",X"FF86",X"FE6F",X"FCD2",X"FA99",X"FAA9",X"FBBA",X"FCE4",X"FBA7",X"F7D3",X"F3CB",X"F071",X"EEE0",X"EE0F",X"F2C8",X"FE63",X"0955",X"11C3",X"1730",X"1452",X"0CC8",X"01BE",X"F95A",X"F6BB",X"F8E0",X"0107",X"0CDC",X"1157",X"1237",X"0AB3",X"FFED",X"FCC5",X"FC97",X"FE34",X"0118",X"0030",X"FEC1",X"FD2B",X"FAD7",X"FB58",X"FCB2",X"FDC2",X"FC4E",X"F7DA",X"F3CF",X"F089",X"EE68",X"EEAC",X"F519",X"0136",X"0BA3",X"131E",X"16DA",X"134E",X"0B57",X"00B9",X"F99B",X"F839",X"FAAC",X"03C8",X"0E83",X"121A",X"10AE",X"0812",X"FDC8",X"FB39",X"FB0A",X"FD22",X"FFC6",X"FEF9",X"FDC3",X"FC70",X"FA65",X"FAFF",X"FC19",X"FC91",X"FA7F",X"F680",X"F319",X"F0C0",X"EDD4",X"ED45",X"F5B2",X"018C",X"0BB0",X"1465",X"15D0",X"10CE",X"08B4",X"FE52",X"F80F",X"F78E",X"FA36",X"04E3",X"0F7D",X"125E",X"0F3D",X"0663",X"FD4E",X"FAD8",X"FB30",X"FE16",X"FF38",X"FDFA",X"FCE7",X"FB7E",X"FA75",X"FB18",X"FC51",X"FC79",X"F9A6",X"F5BB",X"F2B6",X"EFAD",X"EE09",X"EF5D",X"F7D6",X"0374",X"0D54",X"14B1",X"14C9",X"0EF8",X"0656",X"FD85",X"F849",X"F8FF",X"FD1C",X"0868",X"10D5",X"1200",X"0D6F",X"0477",X"FDC1",X"FC7A",X"FCBD",X"FF73",X"FFB0",X"FDE2",X"FC8F",X"FAFC",X"FAF0",X"FC1A",X"FD32",X"FC87",X"F914",X"F5A5",X"F2A4",X"EFF1",X"EE8D",X"F0BD",X"FA25",X"0572",X"0F85",X"168D",X"147F",X"0DD1",X"046F",X"FBC9",X"F888",X"F98C",X"FDE7",X"0949",X"10CF",X"11F5",X"0C5C",X"02A1",X"FCB4",X"FBC1",X"FC96",X"FFDF",X"FFB6",X"FE2C",X"FCD7",X"FB3B",X"FB96",X"FCEB",X"FD77",X"FC80",X"F8E3",X"F4B1",X"F123",X"EFF5",X"EF4C",X"F333",X"FD6C",X"07D6",X"0FD5",X"14E5",X"1289",X"0C3A",X"0332",X"FC38",X"F9EA",X"FB2E",X"009A",X"0B9D",X"11BD",X"11E6",X"0B5B",X"0223",X"FDB0",X"FCF8",X"FDCC",X"FFF3",X"FF43",X"FE28",X"FD4A",X"FC49",X"FC94",X"FD74",X"FD55",X"FB26",X"F70F",X"F3B5",X"F10A",X"F005",X"EF80",X"F4EB",X"FE65",X"08BF",X"10B7",X"1424",X"10D1",X"0A5F",X"00B0",X"FB12",X"F9DC",X"FB33",X"01AD",X"0BF2",X"10A3",X"104D",X"08F2",X"FFF6",X"FCB5",X"FCBA",X"FE98",X"0047",X"FE88",X"FD49",X"FC02",X"FB4D",X"FC6D",X"FD34",X"FCBE",X"FA43",X"F5A0",X"F2BF",X"F0CC",X"EF79",X"EF17",X"F594",X"FFCC",X"0993",X"0FD0",X"11E0",X"0E36",X"0810",X"FFBA",X"FAF7",X"F9E4",X"FB87",X"0266",X"0BF0",X"0FFE",X"0EB2",X"07B6",X"FF7D",X"FC86",X"FCBE",X"FEC4",X"FFD5",X"FE81",X"FD46",X"FC70",X"FC20",X"FD19",X"FE19",X"FD47",X"FA11",X"F589",X"F254",X"F085",X"EFCD",X"F051",X"F770",X"0160",X"0ACB",X"1179",X"12A3",X"0EDE",X"081E",X"FF49",X"FB13",X"FA85",X"FC6D",X"04D0",X"0D59",X"0FE4",X"0DC6",X"05FA",X"FF43",X"FDE7",X"FD68",X"FF3E",X"FFC7",X"FDF5",X"FD6B",X"FCC4",X"FCD0",X"FE2B",X"FE97",X"FD76",X"FA24",X"F5B2",X"F319",X"F165",X"F0B0",X"F206",X"F8D5",X"0276",X"0B33",X"1043",X"10B2",X"0D45",X"0745",X"FFD8",X"FC11",X"FB93",X"FD76",X"0595",X"0D9E",X"0FFD",X"0CB5",X"0566",X"FF80",X"FDC8",X"FDCE",X"FF8F",X"FF3A",X"FE06",X"FDC3",X"FD04",X"FDB2",X"FE9D",X"FE73",X"FCAB",X"F8E5",X"F52B",X"F2B6",X"F14E",X"F1A3",X"F2CE",X"FA1B",X"03B7",X"0BA1",X"102C",X"0F6E",X"0B1B",X"0567",X"FF7E",X"FD41",X"FD4F",X"FEE6",X"06E0",X"0D4A",X"0E3E",X"0AEC",X"03F7",X"FEE4",X"FE04",X"FDFF",X"FF0D",X"FDF6",X"FCC4",X"FC25",X"FBB8",X"FD50",X"FE8F",X"FE19",X"FC4F",X"F823",X"F4AD",X"F319",X"F217",X"F22C",X"F3E7",X"FAF9",X"03E5",X"0B58",X"0F6D",X"0DF2",X"0A01",X"0500",X"FFD5",X"FE01",X"FDDB",X"FF39",X"05BC",X"0BA1",X"0D0B",X"09DE",X"03CF",X"FF5F",X"FE42",X"FE6B",X"FF6E",X"FE48",X"FCEF",X"FC33",X"FB9A",X"FC64",X"FDBA",X"FD3F",X"FB35",X"F775",X"F40A",X"F2C5",X"F205",X"F15C",X"F424",X"FB35",X"02D6",X"09B5",X"0D73",X"0C6C",X"08E8",X"04DF",X"00F5",X"FF55",X"FF54",X"0162",X"070A",X"0BCA",X"0C62",X"0940",X"0366",X"00A4",X"0066",X"FF8D",X"FF6C",X"FE21",X"FC91",X"FC87",X"FC8F",X"FD8B",X"FEAA",X"FD30",X"FAB8",X"F73C",X"F401",X"F2E4",X"F2B6",X"F2C1",X"F6BF",X"FD5C",X"03CA",X"0980",X"0BFB",X"0B5C",X"08CA",X"051B",X"023F",X"00BC",X"003A",X"0233",X"0759",X"0B48",X"0B70",X"07A6",X"02EB",X"00BE",X"0004",X"FFCA",X"FF73",X"FDE1",X"FCAA",X"FC78",X"FD02",X"FE39",X"FEDA",X"FD70",X"FAE1",X"F74B",X"F4E8",X"F438",X"F409",X"F471",X"F7E0",X"FE6C",X"054C",X"09D4",X"0B7B",X"0A2A",X"0783",X"0551",X"03CD",X"02AF",X"02BB",X"04A9",X"08A6",X"0B3E",X"0A4A",X"070D",X"0371",X"01EB",X"0106",X"FFF3",X"FEE4",X"FD2D",X"FC2A",X"FBD0",X"FC3C",X"FD7C",X"FD90",X"FC01",X"F975",X"F608",X"F41D",X"F3A4",X"F391",X"F478",X"F890",X"FEA6",X"05A6",X"0974",X"0A09",X"08FC",X"0636",X"0468",X"0386",X"02B7",X"038B",X"048E",X"0710",X"087C",X"06C3",X"04AA",X"023F",X"0092",X"FFD0",X"FDF4",X"FCC7",X"FBE4",X"FB4C",X"FBCA",X"FCA6",X"FD03",X"FC0C",X"FA20",X"F80E",X"F548",X"F426",X"F497",X"F47E",X"F615",X"FA95",X"0030",X"0611",X"0816",X"082A",X"077D",X"0600",X"055B",X"0558",X"0551",X"0619",X"0682",X"06E0",X"06E8",X"053E",X"040E",X"034F",X"01CF",X"0093",X"FF33",X"FDC6",X"FCC0",X"FBF1",X"FC1F",X"FC5E",X"FBE6",X"FB2B",X"F98F",X"F745",X"F5CB",X"F4AB",X"F46F",X"F572",X"F8CA",X"FDFB",X"035A",X"068C",X"07DC",X"07E1",X"0730",X"06A9",X"05F4",X"0596",X"0570",X"0612",X"06A8",X"069B",X"05C8",X"049D",X"0350",X"0207",X"0099",X"FF3D",X"FDC9",X"FCD7",X"FC19",X"FC2C",X"FC9F",X"FC75",X"FBF2",X"FAFB",X"F93A",X"F775",X"F626",X"F5DF",X"F636",X"F812",X"FC71",X"013E",X"057B",X"07C1",X"078D",X"06C8",X"05CF",X"05B4",X"0647",X"06CC",X"067B",X"0597",X"04CA",X"04B7",X"0483",X"0420",X"02D0",X"0147",X"FF73",X"FE38",X"FD8C",X"FD31",X"FD2E",X"FD52",X"FCC0",X"FBDF",X"FB45",X"FA53",X"F8D9",X"F6EB",X"F63B",X"F676",X"F839",X"FC2D",X"0089",X"03FE",X"0655",X"073B",X"0731",X"06AD",X"06AF",X"06BC",X"06C7",X"0637",X"0528",X"04A1",X"0468",X"044E",X"042C",X"02EE",X"015E",X"FF8A",X"FDEF",X"FD49",X"FCC7",X"FC52",X"FC54",X"FC27",X"FB9A",X"FADA",X"F9D4",X"F859",X"F704",X"F659",X"F654",X"F7C6",X"FAD8",X"FEDC",X"029B",X"04A5",X"0578",X"05CF",X"059C",X"0555",X"0564",X"05BD",X"057C",X"04AD",X"03EC",X"0379",X"0357",X"030C",X"0292",X"01AF",X"FFE2",X"FE72",X"FDCC",X"FD99",X"FD8D",X"FD61",X"FCC5",X"FC05",X"FB9F",X"FB4D",X"FA46",X"F92F",X"F7E4",X"F6F9",X"F751",X"F986",X"FD37",X"012E",X"03C5",X"056E",X"065E",X"065A",X"05F2",X"05E5",X"05BF",X"0551",X"0463",X"03EE",X"0394",X"038D",X"036F",X"02F4",X"01E1",X"0074",X"FEEA",X"FE22",X"FD93",X"FD27",X"FCBD",X"FC38",X"FBA0",X"FB97",X"FB53",X"FA97",X"F994",X"F8AA",X"F80F",X"F871",X"FA2B",X"FD0C",X"0074",X"02EF",X"04A5",X"05F9",X"0686",X"06D0",X"06EC",X"073C",X"0719",X"05F7",X"0488",X"03AA",X"0379",X"03B6",X"0351",X"029C",X"013E",X"FFA4",X"FE80",X"FDEC",X"FD8C",X"FD38",X"FCAD",X"FBFB",X"FB33",X"FAF3",X"FADD",X"FA2B",X"F913",X"F841",X"F809",X"F960",X"FCA3",X"FFF8",X"022D",X"03A0",X"049F",X"0517",X"05BA",X"0689",X"0733",X"0736",X"0646",X"0500",X"0404",X"0397",X"03B1",X"0388",X"029C",X"0174",X"0043",X"FF48",X"FECE",X"FE8B",X"FDE8",X"FD32",X"FC22",X"FB04",X"FA9B",X"FAB5",X"FA4E",X"F9A9",X"F90E",X"F88D",X"F936",X"FB40",X"FE12",X"0093",X"0268",X"0374",X"03F6",X"0494",X"0507",X"05BA",X"0653",X"0605",X"0527",X"0411",X"034A",X"02FD",X"02D0",X"0268",X"0174",X"002D",X"FF33",X"FEBB",X"FEB4",X"FE76",X"FDB5",X"FC85",X"FB5E",X"FAAC",X"FA8B",X"FA3C",X"F9E1",X"F99C",X"F922",X"F8F7",X"FA99",X"FD86",X"0044",X"01D5",X"02B8",X"0370",X"042D",X"050C",X"05D0",X"0645",X"0611",X"051E",X"03ED",X"02E1",X"02B1",X"02C8",X"028D",X"0196",X"002D",X"FF4F",X"FECB",X"FE79",X"FE45",X"FD98",X"FC9C",X"FB97",X"FB09",X"FAB4",X"FA79",X"FA6E",X"FA18",X"F97D",X"F982",X"FA51",X"FC70",X"FF0D",X"0126",X"0231",X"02EF",X"03A8",X"049C",X"0585",X"065A",X"06B3",X"0647",X"0554",X"0456",X"03B9",X"0362",X"02F3",X"0206",X"00B1",X"FFAB",X"FF2D",X"FEFC",X"FEDC",X"FEA6",X"FDFF",X"FCE1",X"FBEF",X"FB75",X"FB01",X"FAC3",X"FAC3",X"FAB9",X"FAA2",X"FAB7",X"FC0A",X"FDF5",X"FFB9",X"00E7",X"01CE",X"02B5",X"035F",X"0416",X"04E3",X"0553",X"0568",X"0535",X"04BA",X"03E6",X"031A",X"02E0",X"02C0",X"0226",X"0162",X"0082",X"0011",X"FFC1",X"FF70",X"FEEA",X"FE19",X"FD60",X"FCE0",X"FC8B",X"FC6D",X"FC79",X"FC2E",X"FBEA",X"FB85",X"FB81",X"FCA1",X"FE6E",X"001D",X"0137",X"01C7",X"02A9",X"0387",X"043E",X"050B",X"0586",X"054E",X"04A7",X"040B",X"036D",X"032B",X"02E6",X"026C",X"0157",X"0031",X"FF59",X"FEB5",X"FE7B",X"FE51",X"FDE6",X"FD2E",X"FC4D",X"FBD5",X"FBA5",X"FBB1",X"FBC0",X"FB87",X"FB2C",X"FB53",X"FBC4",X"FCC1",X"FE24",X"FFD3",X"00F5",X"01B4",X"0227",X"02E0",X"03DC",X"047A",X"04D8",X"0511",X"049D",X"040A",X"034E",X"02C6",X"0284",X"022F",X"019C",X"00C8",X"FFD3",X"FF03",X"FE7D",X"FE59",X"FDFA",X"FD64",X"FC8B",X"FC0C",X"FBC8",X"FBCB",X"FC18",X"FC4C",X"FC32",X"FC68",X"FCC2",X"FD4C",X"FE55",X"FF81",X"00AC",X"018F",X"0232",X"02A4",X"02EE",X"038D",X"0421",X"048F",X"0478",X"03EA",X"0327",X"0266",X"01BD",X"013B",X"009B",X"FFDF",X"FF1C",X"FE7F",X"FDCD",X"FD89",X"FD50",X"FCCA",X"FC67",X"FC02",X"FBC5",X"FB80",X"FB80",X"FB86",X"FBAD",X"FC12",X"FC99",X"FD1B",X"FDEE",X"FF26",X"008C",X"01C4",X"02C0",X"039D",X"0447",X"048B",X"04CA",X"04F5",X"050C",X"04C9",X"043E",X"039B",X"02ED",X"025F",X"0201",X"0152",X"009E",X"FFE1",X"FF2A",X"FEDF",X"FE68",X"FDDD",X"FD79",X"FD15",X"FCF6",X"FCB0",X"FC96",X"FC85",X"FCDC",X"FD30",X"FD6F",X"FDA4",X"FE3C",X"FF80",X"009D",X"0135",X"0205",X"02A6",X"0330",X"0377",X"03E1",X"0419",X"03E8",X"0382",X"02E4",X"0237",X"0190",X"011B",X"00C9",X"0064",X"FFD5",X"FF4A",X"FEBE",X"FE49",X"FDF4",X"FDBC",X"FD88",X"FD50",X"FD42",X"FD0D",X"FCEF",X"FD0A",X"FD54",X"FD9F",X"FDF7",X"FE4D",X"FEBF",X"FFB9",X"0085",X"0137",X"01DE",X"02A3",X"0301",X"0303",X"033B",X"037A",X"038C",X"0382",X"0318",X"027A",X"01C5",X"0112",X"009E",X"0063",X"000A",X"FF9B",X"FF09",X"FE74",X"FDE6",X"FD59",X"FCFA",X"FCF4",X"FCDE",X"FCD2",X"FCAF",X"FCB2",X"FD04",X"FD16",X"FD5B",X"FDC9",X"FE52",X"FEF9",X"FF55",X"0012",X"00C8",X"01CA",X"025E",X"0234",X"023C",X"024D",X"02F2",X"031A",X"02C3",X"0281",X"020A",X"01EB",X"0113",X"0064",X"FF9C",X"FF4C",X"FF4B",X"FF24",X"FE8F",X"FE02",X"FDAD",X"FD2D",X"FCEF",X"FD05",X"FCEE",X"FD1B",X"FD95",X"FDE0",X"FDC2",X"FE03",X"FEA3",X"FF44",X"FF65",X"0006",X"004D",X"00C5",X"018B",X"021D",X"0247",X"021B",X"0225",X"024F",X"0267",X"0279",X"022B",X"0200",X"01C9",X"014B",X"00CD",X"0056",X"0009",X"FFAA",X"FF77",X"FF4C",X"FEEE",X"FE66",X"FE5B",X"FE20",X"FDFB",X"FDE6",X"FDFC",X"FE08",X"FE3D",X"FE78",X"FECA",X"FF77",X"0025",X"0086",X"00F5",X"0181",X"024D",X"02A0",X"031F",X"0369",X"0335",X"0303",X"02E0",X"0276",X"01E3",X"0148",X"00E8",X"00ED",X"0134",X"0111",X"00A6",X"003A",X"FFC1",X"FF0C",X"FEBE",X"FEC9",X"FE9D",X"FE53",X"FE11",X"FDFE",X"FE14",X"FE28",X"FDFB",X"FE30",X"FE7E",X"FEC7",X"FF0F",X"FF3B",X"FFB9",X"0014",X"0057",X"00A4",X"0117",X"01A9",X"01E6",X"01F9",X"01EF",X"01D1",X"01CB",X"0194",X"015E",X"012F",X"00E6",X"00F0",X"00B2",X"004D",X"0017",X"FF90",X"FF29",X"FEC2",X"FE59",X"FE04",X"FDD3",X"FDF5",X"FE00",X"FE0B",X"FE33",X"FE58",X"FE8C",X"FEC5",X"FF43",X"FF89",X"FFF1",X"0040",X"0093",X"00D6",X"00EC",X"0100",X"0100",X"0111",X"00F6",X"00FF",X"0124",X"00F6",X"007D",X"003A",X"0038",X"003F",X"0012",X"001C",X"FFE8",X"FF79",X"FF0C",X"FEC7",X"FE90",X"FE48",X"FE30",X"FE47",X"FE53",X"FE40",X"FE21",X"FE28",X"FE06",X"FDFF",X"FE68",X"FECB",X"FF0C",X"FF7B",X"FFC4",X"FFD2",X"FFF1",X"0022",X"0066",X"009B",X"009C",X"00A2",X"00A7",X"0066",X"004E",X"0043",X"0031",X"003D",X"0032",X"0011",X"000A",X"FFD6",X"FFAA",X"FFA1",X"FF94",X"FF6A",X"FF42",X"FF4B",X"FF3F",X"FF50",X"FF42",X"FF82",X"FF9C",X"FF9B",X"FFBE",X"FFED",X"0021",X"0021",X"0016",X"0050",X"009A",X"00D8",X"0103",X"0159",X"0181",X"0199",X"019D",X"016D",X"0162",X"016E",X"0160",X"0138",X"010D",X"00E8",X"00E2",X"00BA",X"0095",X"0055",X"0046",X"0035",X"001F",X"FFFA",X"FFC3",X"FFC7",X"FFD0",X"FFCE",X"FFD9",X"FFCE",X"FFBE",X"FF72",X"FF5C",X"FF7E",X"FF97",X"FFE1",X"0027",X"0066",X"0067",X"004F",X"0049",X"0034",X"0047",X"005A",X"006C",X"0071",X"0071",X"0072",X"0077",X"0051",X"000B",X"0013",X"0019",X"FFFF",X"FFDE",X"FF7D",X"FF41",X"FF3F",X"FF0B",X"FEDF",X"FECD",X"FF03",X"FF39",X"FF52",X"FF5E",X"FF47",X"FF1B",X"FF19",X"FF1A",X"FF44",X"FF8E",X"FF7A",X"FF98",X"FFD2",X"FFFE",X"0011",X"0059",X"0089",X"00A1",X"00A6",X"0070",X"0035",X"004B",X"0053",X"004D",X"005A",X"0042",X"0054",X"0058",X"0035",X"FFF5",X"FFAB",X"FF8D",X"FF64",X"FF35",X"FF27",X"FF08",X"FED5",X"FEF0",X"FF1D",X"FF4D",X"FF4B",X"FF94",X"FFD2",X"FFC6",X"FFC5",X"FFFD",X"0003",X"0012",X"004A",X"0064",X"0066",X"0084",X"007A",X"0068",X"005F",X"0070",X"0044",X"FFFC",X"0016",X"002E",X"FFF6",X"FFB7",X"FF88",X"FF92",X"FFAE",X"FFC5",X"FFC4",X"FFE4",X"FFCF",X"FFA7",X"FF7D",X"FF76",X"FF8E",X"FF66",X"FF74",X"FF91",X"FFA6",X"FF9E",X"FFBF",X"FFFD",X"002C",X"0031",X"0003",X"0008",X"0024",X"0034",X"004B",X"0041",X"0045",X"003C",X"0065",X"00A6",X"00BA",X"00AA",X"00A7",X"00A5",X"00A2",X"0088",X"004B",X"002A",X"0024",X"0015",X"0015",X"0036",X"0061",X"0030",X"001B",X"0020",X"FFF5",X"FFE8",X"FFFB",X"FFFC",X"0044",X"005E",X"005A",X"004A",X"0068",X"0088",X"00A2",X"00A7",X"0091",X"0074",X"002C",X"0009",X"002F",X"0043",X"0048",X"0016",X"0031",X"003B",X"0024",X"0012",X"FFF6",X"FFE0",X"FFE0",X"FF9E",X"FF70",X"FF76",X"FF85",X"FF65",X"FF6F",X"FF63",X"FF6A",X"FFAB",X"FFEA",X"FFD3",X"FFBA",X"FFCB",X"FFE8",X"FFFF",X"000A",X"FFFC",X"000E",X"000B",X"0035",X"006F",X"0090",X"007D",X"004B",X"003D",X"004F",X"0029",X"001E",X"0017",X"0012",X"0019",X"005C",X"0051",X"0022",X"0022",X"0009",X"FFF1",X"FFF4",X"FFED",X"FFBB",X"FFA1",X"FF84",X"FF64",X"FF38",X"FF3C",X"FF07",X"FEFF",X"FF34",X"FF48",X"FF5B",X"FF99",X"FFB9",X"0002",X"0026",X"0050",X"0049",X"004A",X"FFE8",X"FF7F",X"FF6C",X"FF84",X"FF8C",X"FF9A",X"FF3D",X"FF25",X"FF1D",X"FF42",X"FF33",X"FF0E",X"FF0E",X"FF0F",X"FF06",X"FEF5",X"FEBF",X"FEBF",X"FEC7",X"FEB4",X"FEDA",X"FF32",X"FF71",X"FF85",X"FF7A",X"FF7A",X"FF8F",X"FFB1",X"FFC7",X"FFF9",X"0016",X"0036",X"007B",X"00AD",X"009F",X"009C",X"00B2",X"00B3",X"0093",X"006A",X"006F",X"0072",X"0082",X"00AA",X"008E",X"007B",X"009B",X"00DA",X"00EB",X"00E9",X"00D3",X"0099",X"0062",X"0052",X"004D",X"0036",X"000F",X"0034",X"003C",X"0046",X"005B",X"005C",X"006F",X"0097",X"00CA",X"00E7",X"00DE",X"00B3",X"0083",X"009B",X"0095",X"0081",X"007C",X"0065",X"0058",X"006B",X"0055",X"0028",X"0001",X"FFB5",X"FF6D",X"FF76",X"FF7D",X"FF6F",X"FF9C",X"FFE2",X"FFED",X"FFEB",X"FFEA",X"FFF0",X"FFEC",X"0006",X"002F",X"0027",X"0025",X"0012",X"0011",X"002D",X"0029",X"0014",X"0019",X"0011",X"0057",X"006C",X"006F",X"0066",X"003F",X"000D",X"FFE2",X"FFB5",X"FFCA",X"FFDC",X"0000",X"0010",X"000A",X"0009",X"001B",X"0012",X"FFF2",X"FFED",X"FFB9",X"FFA1",X"FF9C",X"FFAA",X"FFA4",X"FF96",X"FF74",X"FF81",X"FF91",X"FF97",X"FF9F",X"FF8B",X"FF7E",X"FF93",X"FF7C",X"FF56",X"FF68",X"FFAE",X"FFC9",X"FFBB",X"FFA5",X"FFA1",X"FFC4",X"FFBF",X"FF91",X"FF5A",X"FF7F",X"FFC0",X"FFF3",X"FFED",X"FFC5",X"FFB3",X"FFC3",X"FFBE",X"FF93",X"FFB9",X"FFDE",X"FFF0",X"FFE9",X"FFCF",X"FFC4",X"FFCA",X"FFAD",X"FFAC",X"FFF2",X"FFF4",X"FFE0",X"FFE5",X"FFE7",X"FFBB",X"FF96",X"FFA8",X"FFB1",X"FFBC",X"FFA0",X"FF84",X"FF97",X"FFA3",X"FFAB",X"FFA8",X"FFBA",X"FFC1",X"FFBE",X"FFE1",X"FFFD",X"001B",X"001F",X"0041",X"0057",X"002C",X"001F",X"0023",X"0040",X"0078",X"0097",X"009F",X"00C6",X"00C1",X"00BA",X"00A2",X"0090",X"00B3",X"00B2",X"008C",X"004E",X"0057",X"00A7",X"00AC",X"0095",X"003F",X"0012",X"FFF0",X"FFEE",X"000B",X"001F",X"0019",X"FFEB",X"FFC7",X"FFB7",X"FF83",X"FFA1",X"FFF9",X"0017",X"0036",X"0022",X"FFFD",X"FFF1",X"FFA3",X"FF81",X"FF8A",X"FFB1",X"FFC0",X"FFF7",X"0004",X"FFEF",X"FFD0",X"FFAA",X"FF8C",X"FFAE",X"FFD1",X"0007",X"0010",X"001E",X"001D",X"FFD2",X"FFD0",X"000F",X"0039",X"002F",X"002C",X"002F",X"0001",X"0005",X"0001",X"FFF0",X"FFFE",X"0016",X"0068",X"0096",X"009E",X"0086",X"0090",X"0077",X"0068",X"006B",X"0058",X"0043",X"004C",X"003A",X"003D",X"0035",X"003B",X"003C",X"0034",X"0048",X"0018",X"FFCF",X"FFE1",X"0009",X"001A",X"FFF4",X"FFB8",X"FFBA",X"FFB0",X"FF93",X"FFA9",X"FFCA",X"FFBC",X"FFA0",X"FF87",X"FF73",X"FFC0",X"FFC1",X"FFC4",X"FFB5",X"FFAF",X"FFAE",X"FFC2",X"FFC8",X"FFBB",X"FFA6",X"FF90",X"FFA8",X"FFA9",X"FFC1",X"FF9B",X"FF76",X"FF68",X"FF2B",X"FF38",X"FF29",X"FEFB",X"FF31",X"FF9A",X"FFC0",X"FFCE",X"FF84",X"FF53",X"FF6D",X"FF55",X"FF71",X"FF5B",X"FF78",X"FF86",X"FF5A",X"FF61",X"FF81",X"FFAD",X"FFAD",X"FFD9",X"0012",X"0002",X"FFE0",X"FFC9",X"0005",X"0034",X"0014",X"0007",X"0038",X"004F",X"0069",X"008A",X"00B9",X"00B9",X"00C3",X"0099",X"0072",X"0087",X"0080",X"0084",X"0073",X"0051",X"005A",X"003F",X"0031",X"0010",X"0008",X"0031",X"0053",X"0039",X"FFFA",X"FFB8",X"FF9D",X"FFE9",X"001F",X"FFFD",X"FFE7",X"002A",X"0059",X"0061",X"005F",X"0042",X"003F",X"002F",X"000C",X"0019",X"0057",X"00A6",X"00C0",X"00B5",X"00B1",X"00C4",X"00D1",X"00B7",X"009A",X"008B",X"0099",X"00BA",X"00E6",X"00C3",X"0077",X"002B",X"0039",X"0076",X"0084",X"0064",X"0024",X"0025",X"003D",X"0001",X"FFE4",X"FFB3",X"FFB0",X"FFB9",X"FFD1",X"FFE2",X"FFF3",X"FFF5",X"FFCD",X"FFAD",X"FF82",X"FF46",X"FF2B",X"FF21",X"FF5B",X"FF89",X"FF89",X"FFDE",X"FFF1",X"FFF5",X"FFFE",X"FFFF",X"001F",X"005E",X"009E",X"00B1",X"004C",X"FFFC",X"0006",X"000D",X"FFFC",X"FFDF",X"FFC9",X"FFC4",X"FFC7",X"FFBE",X"FFAE",X"FF70",X"FF3F",X"FF69",X"FF8A",X"FF64",X"FF22",X"FEF4",X"FEDE",X"FF04",X"FF1D",X"FF0A",X"FF2C",X"FF3F",X"FF6A",X"FF73",X"FFB3",X"FFE5",X"FFD0",X"FF94",X"FF53",X"FF2B",X"FF27",X"FF59",X"FF89",X"FF66",X"FF5E",X"FF79",X"FFA6",X"FFB7",X"FF97",X"FFA7",X"FF96",X"FFAD",X"FFB0",X"FFC1",X"FFD1",X"FFEE",X"0008",X"0008",X"0002",X"0007",X"000A",X"0035",X"0046",X"002D",X"0031",X"000D",X"0005",X"000A",X"FFCC",X"FFB4",X"FFE6",X"003A",X"00AA",X"00A1",X"0091",X"008E",X"008B",X"0079",X"0069",X"004F",X"005A",X"006F",X"0053",X"004A",X"003D",X"0033",X"0009",X"0018",X"0038",X"0062",X"0064",X"0039",X"FFF5",X"FFDD",X"FFC2",X"FFE1",X"001D",X"0045",X"0021",X"FFFD",X"FFCC",X"FFAF",X"FFD5",X"FFEF",X"0015",X"0041",X"0042",X"005D",X"004E",X"0035",X"0060",X"007E",X"009F",X"00B7",X"00C1",X"0093",X"0076",X"0072",X"004F",X"0032",X"0002",X"0017",X"001A",X"0012",X"001A",X"001B",X"000A",X"FFE5",X"FFE6",X"FFEB",X"FFDD",X"FFD1",X"FFD4",X"0009",X"001C",X"FFF6",X"FFE4",X"FFDF",X"0000",X"001C",X"003A",X"0070",X"0079",X"0057",X"0062",X"0038",X"000E",X"0015",X"0012",X"0015",X"003A",X"0054",X"004D",X"003E",X"0026",X"0012",X"FFFF",X"FFF8",X"FFEE",X"FFEC",X"FFCD",X"FFC3",X"FFBD",X"FFA1",X"FF95",X"FFA0",X"FF6E",X"FF48",X"FF41",X"FF6B",X"FF83",X"FF6C",X"FF60",X"FF85",X"FFAC",X"FF9F",X"FF8C",X"FF78",X"FF90",X"FFBF",X"FFB0",X"FF9F",X"FF6B",X"FF32",X"FF48",X"FF55",X"FF6B",X"FFB2",X"FFF9",X"0003",X"0026",X"002C",X"FFFB",X"FFAE",X"FFA2",X"FFC6",X"FFFF",X"003B",X"0010",X"FFD1",X"FFEA",X"FFF2",X"FFED",X"FFCB",X"FFB4",X"FFC9",X"FFBD",X"FF94",X"FF75",X"FF77",X"FF84",X"FFC0",X"FFE1",X"0004",X"0017",X"0018",X"0026",X"0027",X"FFF8",X"000C",X"0017",X"0031",X"005A",X"0055",X"0055",X"0058",X"003C",X"0028",X"FFFF",X"0018",X"0042",X"0045",X"001A",X"003D",X"0074",X"005C",X"0039",X"0020",X"0027",X"002B",X"001A",X"0030",X"002D",X"0029",X"0010",X"0013",X"0017",X"0039",X"0042",X"002E",X"FFFF",X"0006",X"000A",X"FFEB",X"FFF3",X"FFF0",X"FFFF",X"000A",X"0028",X"0052",X"00A7",X"0093",X"0053",X"004E",X"0054",X"004D",X"003C",X"003D",X"0040",X"0015",X"001E",X"0023",X"002E",X"0034",X"000F",X"FFD3",X"FFCA",X"FFEE",X"FFF2",X"0002",X"FFF3",X"FFD3",X"FFE1",X"FFE6",X"0009",X"0019",X"0053",X"0065",X"004F",X"005A",X"004F",X"0048",X"004A",X"0029",X"0056",X"0045",X"003F",X"0053",X"0077",X"0075",X"002C",X"FFF7",X"0029",X"0056",X"005F",X"FFFF",X"FFAF",X"FFB5",X"FFAF",X"FF8C",X"FF5C",X"FF57",X"FF5F",X"FF42",X"FF17",X"FF03",X"FEE7",X"FEF0",X"FEEC",X"FEF9",X"FF32",X"FF2E",X"FF35",X"FF31",X"FF1F",X"FF12",X"FF0E",X"FF09",X"FEEF",X"FEF9",X"FF2C",X"FF4A",X"FF4E",X"FF79",X"FF9C",X"FFAA",X"FFA9",X"FF90",X"FF87",X"FF9A",X"FF90",X"FF88",X"FF7E",X"FF81",X"FF77",X"FF75",X"FF6A",X"FF7E",X"FFAF",X"FFEE",X"FFFA",X"0001",X"002E",X"0030",X"0000",X"000B",X"000A",X"FFF0",X"000E",X"003B",X"0056",X"0066",X"0055",X"0008",X"0008",X"001D",X"004A",X"0074",X"0063",X"0066",X"004C",X"0057",X"0042",X"0030",X"0015",X"0013",X"002F",X"002D",X"0031",X"0059",X"0048",X"0016",X"FFEB",X"FFDD",X"0002",X"000B",X"0024",X"006C",X"0062",X"003B",X"003D",X"0037",X"0056",X"0066",X"0079",X"0092",X"009D",X"0052",X"001A",X"0007",X"FFF6",X"FFE8",X"FFE8",X"FFD5",X"FFF7",X"000D",X"0002",X"FFE9",X"FFEF",X"FFCA",X"FFCA",X"FFD8",X"FFFD",X"FFFF",X"0017",X"FFFD",X"FFFC",X"000D",X"000C",X"0003",X"FFFE",X"0009",X"0039",X"0054",X"0072",X"004F",X"0026",X"0029",X"003C",X"003D",X"0027",X"0049",X"00AE",X"00D8",X"00CB",X"008F",X"0071",X"0050",X"003C",X"0047",X"0045",X"001F",X"000B",X"0001",X"0001",X"001B",X"0012",X"FFFE",X"FFD6",X"FFDB",X"FFD8",X"FFEC",X"0028",X"0016",X"0005",X"FFFA",X"FFEC",X"FFFA",X"0028",X"002B",X"0024",X"0020",X"0038",X"0010",X"FFD0",X"FFC7",X"FFAC",X"FF89",X"FF98",X"FFB3",X"FFD4",X"FFE2",X"FFCD",X"FFAE",X"FFAA",X"FFA9",X"FFAB",X"FF82",X"FF8B",X"FF8A",X"FF95",X"FF99",X"FF5E",X"FF4E",X"FF5D",X"FF84",X"FF6A",X"FF66",X"FF66",X"FF55",X"FF65",X"FF64",X"FF79",X"FF9A",X"FF9E",X"FF84",X"FFC8",X"FFF3",X"0006",X"0027",X"0047",X"001F",X"0002",X"0001",X"0004",X"FFFC",X"FFEC",X"FFD1",X"0003",X"0017",X"0004",X"FFFB",X"FFEF",X"FFDB",X"FFE2",X"FFEA",X"000F",X"0005",X"FFFF",X"FFF8",X"FFFF",X"0002",X"000F",X"000A",X"0043",X"0059",X"0061",X"0046",X"0032",X"0027",X"0011",X"0005",X"FFDF",X"FFCC",X"FFEA",X"0003",X"0003",X"FFEE",X"FFFD",X"FFF0",X"FFE2",X"FFC7",X"FFB3",X"FFAB",X"FFF4",X"002C",X"0009",X"FFB8",X"FFBA",X"FFC8",X"FFC4",X"FFF0",X"FFE6",X"FFD7",X"001C",X"002E",X"0001",X"000F",X"003D",X"0024",X"004D",X"0052",X"003A",X"0032",X"0043",X"004D",X"0073",X"007B",X"0061",X"004B",X"001D",X"002F",X"0059",X"0068",X"0061",X"0051",X"003A",X"0014",X"0009",X"0018",X"0021",X"0024",X"0024",X"0034",X"002D",X"0026",X"FFFB",X"FFF3",X"0001",X"FFFA",X"FFE7",X"FFC3",X"FFA2",X"FFAF",X"FFE0",X"FFE5",X"0009",X"003D",X"0038",X"FFF5",X"FFF1",X"FFFD",X"0009",X"0034",X"001B",X"0003",X"0020",X"0005",X"0003",X"FFEE",X"FFD5",X"FFE3",X"FF95",X"FF5A",X"FF42",X"FF53",X"FF85",X"FFA2",X"FF9C",X"FFA9",X"FF9B",X"FFCB",X"FFF8",X"0010",X"0002",X"FFEC",X"FFF8",X"FFD7",X"FFA7",X"FF81",X"FF83",X"FF61",X"FF21",X"FF3B",X"FF4D",X"FF20",X"FF1C",X"FF18",X"FF20",X"FF4E",X"FF56",X"FF79",X"FF84",X"FF64",X"FF86",X"FFAB",X"FFB0",X"FF93",X"FF99",X"FFBB",X"FFF9",X"0006",X"0023",X"0076",X"0064",X"0074",X"008B",X"005F",X"0075",X"0079",X"006C",X"0053",X"0050",X"0041",X"0005",X"FFF2",X"FFF0",X"FFFF",X"0012",X"003C",X"003E",X"0035",X"0041",X"003B",X"0038",X"0042",X"006C",X"0071",X"007B",X"0065",X"0044",X"0017",X"FFF7",X"FFD4",X"FFE6",X"0021",X"0006",X"FFD3",X"FFD2",X"FFF6",X"001E",X"0030",X"0016",X"FFF1",X"FFEA",X"FFE0",X"FFD3",X"FFBB",X"FFC0",X"FFDA",X"FFD3",X"FFDA",X"FFE2",X"FFED",X"FFFD",X"0015",X"0044",X"0066",X"0030",X"0033",X"0034",X"000B",X"FFFC",X"FFF2",X"FFF6",X"0022",X"0029",X"0041",X"005D",X"0077",X"0083",X"0082",X"007C",X"0092",X"0075",X"0091",X"0099",X"00A2",X"009E",X"008D",X"007C",X"005E",X"0039",X"002D",X"0041",X"0018",X"0020",X"0023",X"FFE0",X"FFB8",X"FFE5",X"FFF6",X"FFFA",X"0013",X"FFFD",X"FFF7",X"FFFC",X"000A",X"FFFD",X"001E",X"0025",X"0002",X"FFF6",X"FFDC",X"FFB7",X"FF9E",X"FFAE",X"FFC8",X"FFCA",X"FFA8",X"FFA0",X"FF83",X"FF4B",X"FF52",X"FF50",X"FF34",X"FF24",X"FF63",X"FF58",X"FF6D",X"FFBC",X"FFAE",X"FF9F",X"FFBE",X"FFB4",X"FFBF",X"FFD7",X"FFA6",X"FF9A",X"FFCA",X"FF9C",X"FF9E",X"FFD1",X"FFA2",X"FF9E",X"FFA2",X"FFAA",X"FFAF",X"FF96",X"FFB6",X"FF8C",X"FF73",X"FF65",X"FF75",X"FF81",X"FF72",X"FFB2",X"FFFA",X"FFF9",X"FFC8",X"FFBE",X"FFA5",X"FFAC",X"FFBE",X"FFA9",X"FF81",X"FFB8",X"FFDE",X"FFEF",X"FFBF",X"FFBD",X"FFDC",X"FFFF",X"FFFE",X"000A",X"0014",X"0032",X"000A",X"0006",X"0048",X"007D",X"007F",X"0071",X"0080",X"00A0",X"00AC",X"00B1",X"00B9",X"0092",X"004C",X"001F",X"0027",X"002B",X"002B",X"0017",X"0001",X"FFE9",X"FFEF",X"FFE0",X"FFEC",X"FFED",X"FFDD",X"FFFF",X"0032",X"0030",X"0036",X"0029",X"FFF5",X"FFD0",X"000A",X"0002",X"FFF7",X"FFE4",X"FFE4",X"FFDD",X"FFDA",X"FFE4",X"FFEB",X"FFEB",X"FFF6",X"002A",X"0051",X"0056",X"0053",X"0069",X"005E",X"0044",X"0036",X"000A",X"FFE7",X"FFEA",X"FFB6",X"FFB3",X"FFD2",X"FFE2",X"FFF0",X"002D",X"0032",X"0019",X"FFF9",X"000E",X"0039",X"000F",X"001B",X"003B",X"0005",X"FFF1",X"FFFE",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000");
	--constant sound2 : table_type := (X"0005",X"0007",X"0004",X"000E",X"001A",X"004A",X"0067",X"0034",X"0031",X"006E",X"00A0",X"009D",X"0072",X"0054",X"003A",X"003E",X"0031",X"0033",X"0053",X"0075",X"0062",X"0068",X"008F",X"0098",X"0095",X"0084",X"006B",X"0055",X"0074",X"0084",X"008E",X"004D",X"0005",X"FFD5",X"FFC7",X"FFCE",X"FFA5",X"FF80",X"FF5F",X"FF78",X"FF89",X"FF77",X"FF97",X"FF86",X"FF78",X"FFB0",X"FFD7",X"FFD7",X"FFEC",X"FFF3",X"FFE6",X"FFDD",X"FFF6",X"FFD3",X"FFB9",X"FFA0",X"FF7A",X"FF6F",X"FF39",X"FF2B",X"FF29",X"FF37",X"FF4C",X"FF81",X"FFD5",X"0001",X"0033",X"006A",X"0021",X"FFDE",X"FFD7",X"FFEE",X"0006",X"0003",X"0013",X"FFF8",X"FFD4",X"FFF3",X"FFDD",X"FFC4",X"FFCB",X"FFF3",X"000E",X"0027",X"002B",X"0020",X"000E",X"FFF7",X"FFF6",X"FFF3",X"FFF9",X"0011",X"001E",X"0011",X"FFE0",X"FFAF",X"FF99",X"FF8B",X"FFAB",X"FFD6",X"FFED",X"FFF7",X"0013",X"000B",X"FFD8",X"FFA0",X"FF8B",X"FF9C",X"FFB2",X"FFD0",X"FFD8",X"FF82",X"FF22",X"FF49",X"FF75",X"FF5E",X"FF3F",X"FF13",X"FEF7",X"FF16",X"FF63",X"FF88",X"FFB6",X"FFAD",X"FFA4",X"FFC9",X"FFB6",X"FFCB",X"FFE5",X"FFEB",X"0001",X"FFE9",X"0009",X"0003",X"FFF6",X"FFFE",X"0010",X"0038",X"0062",X"008F",X"0093",X"008F",X"0094",X"00D5",X"00F3",X"00BE",X"009F",X"00BA",X"00D2",X"00C8",X"00C2",X"009B",X"0077",X"0051",X"0088",X"00BF",X"00AD",X"00A0",X"00CA",X"00C9",X"009B",X"009F",X"009D",X"00B7",X"0089",X"005B",X"0050",X"0012",X"FFE3",X"FFD1",X"FFCB",X"FFAA",X"FFB0",X"FFB6",X"FFA6",X"FF87",X"FFA9",X"FFDA",X"FFEF",X"FFFC",X"FFF6",X"FFE7",X"FFE1",X"FFF7",X"0001",X"0006",X"FFB1",X"FF4A",X"FF2A",X"FF23",X"FF49",X"FF61",X"FF68",X"FF55",X"FF5C",X"FF6D",X"FF69",X"FF89",X"FFD1",X"FFF1",X"FFFE",X"FFD4",X"FFC5",X"FFD4",X"FFAC",X"FF8B",X"FF74",X"FF4D",X"FF6A",X"FF83",X"FF91",X"FF81",X"FF70",X"FF7B",X"FFB3",X"0000",X"0024",X"0054",X"0098",X"009F",X"0098",X"007F",X"005D",X"0039",X"0023",X"0015",X"FFFF",X"FFEA",X"FFC8",X"FF91",X"FF8F",X"FFD1",X"FFE8",X"FFDE",X"000D",X"002E",X"0078",X"00A4",X"00AB",X"006F",X"0024",X"0001",X"FFFB",X"0009",X"FFF0",X"FFBB",X"FFAB",X"FF81",X"FF43",X"FF07",X"FF05",X"FF10",X"FF6B",X"FFD6",X"FFFA",X"FFFD",X"FFFB",X"0002",X"0000",X"FFC8",X"FFA8",X"FFA4",X"FF8C",X"FF7A",X"FFB9",X"FFD8",X"FFB3",X"FFAC",X"FF84",X"FF52",X"FF39",X"FF4E",X"FFA8",X"0008",X"005F",X"0029",X"0006",X"FFBD",X"FFD7",X"0014",X"002A",X"0025",X"0022",X"0027",X"0014",X"0004",X"0014",X"0036",X"004D",X"0044",X"0053",X"0070",X"0094",X"00AA",X"00B1",X"00EC",X"00FE",X"00E3",X"00C9",X"00AA",X"0087",X"0069",X"004C",X"002F",X"0015",X"000C",X"0025",X"0053",X"0094",X"00E9",X"0107",X"00F6",X"00E2",X"00C4",X"00CE",X"00DA",X"00C3",X"009B",X"00B1",X"00BE",X"0078",X"003A",X"000F",X"FFED",X"FFB5",X"FF86",X"FFA6",X"FFCE",X"000B",X"001E",X"0030",X"0050",X"0019",X"FFE5",X"FFC3",X"FFBE",X"FF99",X"FF6C",X"FF40",X"FEF7",X"FEAB",X"FE9E",X"FE9E",X"FEBF",X"FEF5",X"FF64",X"FF48",X"FF39",X"FF6E",X"FFBE",X"FFFA",X"001D",X"002F",X"0010",X"FFFD",X"FFF2",X"FFDE",X"FFC9",X"FFC0",X"FF8E",X"FF33",X"FF3C",X"FF5A",X"0292",X"0152",X"007B",X"01EF",X"00BF",X"00FC",X"007D",X"0040",X"018B",X"003E",X"FDD5",X"FDA9",X"FE09",X"FC72",X"FC5D",X"FCA7",X"FD33",X"FDDA",X"FE46",X"FE24",X"000A",X"013C",X"014F",X"01CC",X"031F",X"02F9",X"034C",X"02A7",X"017A",X"0136",X"0119",X"FF6A",X"FE7A",X"FECC",X"FDFF",X"FCB6",X"FCFE",X"FD7F",X"FE75",X"FFA3",X"007B",X"013B",X"02AF",X"03AC",X"0455",X"0452",X"03AA",X"0322",X"01F5",X"FFEE",X"FDD1",X"FC71",X"FAD8",X"F944",X"F8E2",X"F95F",X"F9CA",X"FB18",X"FD1F",X"FF53",X"0220",X"04EB",X"06E0",X"08B0",X"0A1C",X"09E3",X"0817",X"0519",X"01C8",X"FE8F",X"F9E0",X"F5DF",X"F3E0",X"F295",X"F254",X"F31B",X"F5D9",X"FA29",X"FF08",X"047A",X"0A64",X"0FBA",X"13B8",X"161E",X"15D1",X"126C",X"0B01",X"04ED",X"FEC0",X"F54F",X"ED43",X"E924",X"E6B9",X"E575",X"E75A",X"ECC9",X"F4E8",X"FE56",X"083C",X"11DD",X"1AC8",X"2141",X"2444",X"22BE",X"1C96",X"1240",X"092A",X"FE99",X"F06D",X"E5BE",X"DFBD",X"DB2E",X"D932",X"DC1F",X"E471",X"EF1E",X"FA79",X"06D9",X"12F0",X"1CD2",X"2422",X"27B2",X"25FC",X"1F88",X"14F9",X"0B1A",X"0044",X"F276",X"E742",X"E0F8",X"DC12",X"D83B",X"D9A4",X"E195",X"EBDE",X"F735",X"04DD",X"1268",X"1D86",X"2619",X"2B40",X"2AB6",X"24EE",X"1A11",X"0F5F",X"034C",X"F4DC",X"E7F9",X"DFF6",X"D9F4",X"D54E",X"D59D",X"DB21",X"E534",X"F1C0",X"FFCF",X"0E72",X"1B8C",X"25FB",X"2CDD",X"2E6E",X"2A46",X"2105",X"141E",X"07D6",X"FA4E",X"EB12",X"DFD7",X"D93F",X"D4D5",X"D272",X"D571",X"DF17",X"EB52",X"F914",X"0855",X"1711",X"239B",X"2C93",X"30F9",X"2F69",X"282C",X"1BD6",X"0E12",X"00C4",X"F1AE",X"E365",X"DA7A",X"D533",X"D161",X"D183",X"D799",X"E334",X"F0CC",X"0023",X"1057",X"1E98",X"29BF",X"30DE",X"32F6",X"2E9C",X"24D5",X"16E8",X"08AE",X"FA72",X"EB15",X"DE2A",X"D6BA",X"D299",X"D061",X"D2F3",X"DBC1",X"E88E",X"F82A",X"084C",X"1705",X"2459",X"2E96",X"33F1",X"32D2",X"2C5D",X"20ED",X"11AF",X"0261",X"F313",X"E3B5",X"D818",X"D292",X"D023",X"CFC7",X"D4CA",X"E03B",X"EF4A",X"FFC1",X"0FF8",X"1E64",X"2B2C",X"341E",X"368A",X"31A0",X"2807",X"1B17",X"0AD9",X"FA3E",X"EA9D",X"DC9A",X"D39B",X"CF99",X"CE5C",X"D084",X"D818",X"E63E",X"F712",X"06A6",X"15F4",X"2574",X"313D",X"3633",X"354C",X"2E99",X"22ED",X"13BF",X"0280",X"F27C",X"E3DE",X"D811",X"D15F",X"CEDD",X"CF7F",X"D401",X"DD96",X"ECDB",X"FE08",X"0D9F",X"1C0B",X"29A2",X"333B",X"35FD",X"3257",X"2975",X"1C9C",X"0CCE",X"FC55",X"EC8E",X"DF59",X"D607",X"D196",X"D0AB",X"D267",X"D86A",X"E3C8",X"F399",X"03FC",X"1269",X"1FCF",X"2BF9",X"337C",X"33F4",X"2E51",X"23FE",X"169E",X"06D0",X"F71A",X"E8B4",X"DCF5",X"D570",X"D28D",X"D2B1",X"D538",X"DC1B",X"E881",X"F887",X"07F2",X"151F",X"2218",X"2D85",X"3342",X"31F7",X"2AC8",X"1F86",X"124C",X"0264",X"F29F",X"E537",X"DAB2",X"D4CA",X"D2F0",X"D3AD",X"D6DD",X"DEC4",X"EC84",X"FD04",X"0B2A",X"17F5",X"2563",X"2FAD",X"335C",X"30F5",X"284F",X"1BD1",X"0DFE",X"FDF6",X"EE3A",X"E133",X"D857",X"D3AD",X"D28A",X"D434",X"D8D3",X"E1C9",X"F132",X"0295",X"0FAD",X"1BFA",X"298A",X"32AB",X"3425",X"2F5C",X"24FD",X"17EA",X"09BA",X"F8FE",X"E941",X"DDB1",X"D6BD",X"D341",X"D24E",X"D519",X"DBB6",X"E658",X"F6BF",X"0750",X"1379",X"20DF",X"2E24",X"345E",X"3342",X"2D15",X"21EE",X"13A3",X"03EB",X"F3F8",X"E540",X"DAA2",X"D50B",X"D2C5",X"D2FC",X"D6DF",X"DEB7",X"EB15",X"FC3D",X"0C39",X"1827",X"2593",X"31AD",X"3584",X"3262",X"2A4B",X"1D99",X"0ED6",X"FECE",X"EED1",X"E0F3",X"D7AE",X"D351",X"D210",X"D372",X"D889",X"E1F5",X"F01E",X"0203",X"10A6",X"1BD6",X"2955",X"341F",X"350E",X"2F52",X"25A1",X"189E",X"0982",X"F944",X"E970",X"DCD4",X"D586",X"D2A8",X"D1E5",X"D47D",X"DB10",X"E594",X"F5E3",X"07F6",X"147D",X"1F01",X"2CCF",X"3582",X"33C4",X"2CC9",X"221D",X"1461",X"050F",X"F500",X"E511",X"DA06",X"D4EC",X"D2C5",X"D250",X"D657",X"DEA4",X"EA23",X"FA82",X"0BC0",X"1779",X"2287",X"2FA4",X"35E1",X"3226",X"29B3",X"1E2E",X"0FF5",X"0069",X"F030",X"E194",X"D7F8",X"D424",X"D2F9",X"D37E",X"D893",X"E1FD",X"EEF7",X"FFCE",X"101D",X"1ABF",X"2654",X"3181",X"348F",X"2F0F",X"2572",X"194D",X"0A73",X"FB15",X"EBAA",X"DE6A",X"D60E",X"D415",X"D3BA",X"D52E",X"DB60",X"E5AB",X"F3AF",X"052C",X"13FE",X"1D0E",X"2886",X"330B",X"337D",X"2BBC",X"213A",X"1428",X"0500",X"F5CA",X"E71C",X"DB08",X"D4AC",X"D3EC",X"D4B3",X"D777",X"DEC3",X"E9BD",X"F926",X"0B1A",X"17A8",X"208C",X"2BFA",X"34AC",X"3256",X"28E8",X"1CE2",X"0FAF",X"0127",X"F1C7",X"E2F5",X"D8AD",X"D4F9",X"D4CC",X"D595",X"D9B5",X"E22C",X"EE5A",X"FF94",X"10AE",X"1AD7",X"2482",X"3032",X"34ED",X"3039",X"264C",X"192B",X"0AA7",X"FC7B",X"ED94",X"DEAE",X"D5CA",X"D43B",X"D4B7",X"D5EE",X"DBC7",X"E59C",X"F395",X"05CA",X"150F",X"1DA5",X"2873",X"33D2",X"3506",X"2D02",X"2229",X"14C2",X"0519",X"F665",X"E78D",X"DA0B",X"D354",X"D386",X"D4AD",X"D713",X"DE76",X"E96D",X"F930",X"0BE9",X"18F1",X"2103",X"2C6E",X"3559",X"337C",X"2A0A",X"1D52",X"0EEF",X"FFF7",X"F106",X"E1FD",X"D6B1",X"D281",X"D3A1",X"D551",X"D9CA",X"E240",X"EE9A",X"000B",X"11F9",X"1C8E",X"2564",X"3059",X"3571",X"30DC",X"25EA",X"17B0",X"0884",X"FA6A",X"EC4D",X"DDB4",X"D428",X"D2A7",X"D4BC",X"D76B",X"DCBC",X"E5B4",X"F405",X"0715",X"1673",X"1ECA",X"280F",X"328E",X"34D3",X"2D13",X"2020",X"11E7",X"03E9",X"F652",X"E7F7",X"DA5E",X"D36B",X"D40E",X"D69E",X"D962",X"DF1C",X"E9B9",X"FA83",X"0D9F",X"1988",X"20E8",X"2AE5",X"32F4",X"3242",X"28D9",X"1A22",X"0B10",X"FF0D",X"F258",X"E299",X"D655",X"D33F",X"D592",X"D789",X"DB07",X"E1FD",X"EEC2",X"01C8",X"1327",X"1BB4",X"23CB",X"2F17",X"3447",X"2F37",X"2355",X"1512",X"0725",X"FA83",X"ED3E",X"DE17",X"D482",X"D424",X"D715",X"D90B",X"DD4D",X"E645",X"F5C4",X"09A7",X"17FA",X"1F88",X"2839",X"31B2",X"33D2",X"2B5F",X"1D57",X"0E6A",X"018A",X"F595",X"E6C6",X"D8B2",X"D374",X"D592",X"D811",X"DAF0",X"E0FD",X"ECE2",X"FF28",X"11A9",X"1C93",X"241B",X"2D85",X"33CF",X"3104",X"25A0",X"1667",X"0748",X"FABE",X"EE07",X"DF5E",X"D48C",X"D288",X"D5DD",X"D9BD",X"DE42",X"E650",X"F523",X"0906",X"190D",X"2164",X"2846",X"3049",X"334D",X"2C6C",X"1DC3",X"0CD0",X"FF4E",X"F3E5",X"E601",X"D849",X"D1BA",X"D370",X"D842",X"DCE4",X"E27C",X"ED1A",X"FEF5",X"1277",X"1EC8",X"252F",X"2C4A",X"323A",X"309A",X"2587",X"14CE",X"046E",X"F89B",X"ED8F",X"DF9A",X"D458",X"D21D",X"D6B4",X"DC34",X"E0FA",X"E7E4",X"F598",X"09B8",X"1A5B",X"2283",X"2826",X"2E9E",X"3199",X"2B77",X"1CA8",X"0AE4",X"FD49",X"F327",X"E6FE",X"D9CB",X"D2BE",X"D450",X"D94B",X"DE79",X"E3E1",X"ED4E",X"FE48",X"11A7",X"1E0C",X"2433",X"2A95",X"2FB7",X"2E83",X"249D",X"1448",X"03BF",X"F828",X"EE2E",X"E12A",X"D5EC",X"D311",X"D6B5",X"DBE7",X"E112",X"E7A0",X"F443",X"07B7",X"18CB",X"21A6",X"273A",X"2D5C",X"302C",X"2AB7",X"1D18",X"0BB7",X"FDA5",X"F382",X"E7E8",X"DB24",X"D3D3",X"D467",X"D8EE",X"DE46",X"E415",X"ED91",X"FDF5",X"119D",X"1F21",X"25E3",X"2BD6",X"3087",X"2ECA",X"24A7",X"1490",X"0429",X"F749",X"EC74",X"E042",X"D5D1",X"D23B",X"D553",X"DB17",X"E156",X"E942",X"F678",X"09B9",X"1B1A",X"2505",X"2ADC",X"2F3F",X"30A2",X"2B0C",X"1D24",X"0ABF",X"FB18",X"F020",X"E4FB",X"D90C",X"D1E1",X"D299",X"D814",X"DF3C",X"E6E4",X"F10B",X"01A1",X"152A",X"22A2",X"294A",X"2E44",X"3166",X"2E97",X"23D2",X"1257",X"008B",X"F2F2",X"E83E",X"DCD6",X"D385",X"D103",X"D4B5",X"DBC0",X"E3C3",X"ECAF",X"FA20",X"0D12",X"1E4A",X"27D5",X"2D17",X"308B",X"2FF5",X"286C",X"195C",X"0680",X"F687",X"EB78",X"E0EE",X"D686",X"D110",X"D2BD",X"D8FE",X"E0F1",X"E9A3",X"F4C2",X"059C",X"18AC",X"25D9",X"2BFE",X"2F90",X"30DB",X"2C3B",X"2009",X"0E09",X"FC3B",X"EF0B",X"E4F3",X"DA79",X"D25A",X"D14F",X"D603",X"DD8B",X"E66E",X"F089",X"FEC4",X"11D7",X"2200",X"2A50",X"2EC7",X"30F0",X"2E42",X"251D",X"1587",X"02B9",X"F31F",X"E848",X"DE7C",X"D4CD",X"D07C",X"D357",X"DA74",X"E2C6",X"EC41",X"F8E5",X"0A4E",X"1C4D",X"27E6",X"2DAC",X"305C",X"2FF4",X"29B4",X"1C32",X"09F1",X"F8D5",X"EC49",X"E15B",X"D753",X"D125",X"D0FD",X"D612",X"DE37",X"E7D5",X"F305",X"0292",X"1588",X"2424",X"2BE5",X"3025",X"3134",X"2C9F",X"21B8",X"1193",X"FF70",X"F045",X"E521",X"DB61",X"D33C",X"D086",X"D3F0",X"DAE0",X"E412",X"EEE6",X"FC7C",X"0E41",X"1F7C",X"29FA",X"2F2B",X"31A4",X"2F88",X"271B",X"189A",X"0661",X"F5CA",X"E9B4",X"DF90",X"D65A",X"D164",X"D2D2",X"D8C2",X"E153",X"EB2C",X"F74F",X"07A8",X"19BB",X"269B",X"2D46",X"3116",X"310B",X"2AE8",X"1E6F",X"0D9A",X"FC19",X"ED95",X"E2A9",X"D99A",X"D302",X"D1D6",X"D627",X"DDAF",X"E7A2",X"F31C",X"0153",X"12F9",X"2241",X"2B29",X"2FC2",X"30C4",X"2C79",X"221D",X"12E2",X"00FE",X"F12D",X"E574",X"DC0E",X"D458",X"D170",X"D4A3",X"DB5E",X"E44D",X"EF1F",X"FC83",X"0D86",X"1DE6",X"2894",X"2E58",X"30EA",X"2E53",X"2559",X"17A0",X"0687",X"F5F7",X"E8F9",X"DF2D",X"D709",X"D265",X"D3B2",X"D98A",X"E1A8",X"EBD3",X"F8D9",X"08DB",X"19A7",X"264C",X"2D5C",X"3090",X"2F6D",X"28B0",X"1C19",X"0B97",X"FABF",X"EC6A",X"E16A",X"D8FC",X"D353",X"D287",X"D6F4",X"DEC4",X"E8AC",X"F4F2",X"0436",X"1546",X"230A",X"2BDC",X"3074",X"300A",X"2AA1",X"1F9D",X"0F8F",X"FE5E",X"EF97",X"E3D4",X"DA77",X"D405",X"D20C",X"D580",X"DCB1",X"E5E0",X"F12D",X"005F",X"1248",X"2093",X"29F2",X"2FEE",X"30E6",X"2C1F",X"220F",X"12F2",X"0181",X"F1DB",X"E58A",X"DBA9",X"D482",X"D1D0",X"D414",X"DA8B",X"E450",X"EFB1",X"FDD4",X"0F88",X"1F34",X"2964",X"2FC2",X"319E",X"2D4D",X"237A",X"153E",X"03BB",X"F36A",X"E6A1",X"DC9D",X"D4F0",X"D184",X"D365",X"D992",X"E2EF",X"EEAB",X"FCB5",X"0E03",X"1DFD",X"28DC",X"2FBE",X"31E3",X"2E30",X"252C",X"1703",X"0587",X"F541",X"E7E8",X"DD45",X"D5B5",X"D237",X"D356",X"D8E6",X"E261",X"EEB5",X"FC9A",X"0D54",X"1D49",X"28C0",X"302C",X"3290",X"2EED",X"25CA",X"1857",X"070F",X"F614",X"E811",X"DD38",X"D58C",X"D1F8",X"D311",X"D853",X"E198",X"EDCB",X"FC1E",X"0D3B",X"1CC9",X"27F6",X"2FCC",X"32C6",X"2EF7",X"256B",X"177D",X"061D",X"F5AC",X"E812",X"DC72",X"D458",X"D177",X"D349",X"D8D4",X"E1EF",X"EDE5",X"FC85",X"0E11",X"1DA3",X"281D",X"2F0D",X"322F",X"2EB1",X"24B0",X"1654",X"0554",X"F4E0",X"E74A",X"DC35",X"D42E",X"D137",X"D3A8",X"D9D6",X"E329",X"EF94",X"FE3E",X"0FB1",X"1F64",X"29A1",X"2FF1",X"3243",X"2E40",X"23CA",X"1511",X"039A",X"F33A",X"E60A",X"DB54",X"D3DB",X"D182",X"D48B",X"DB0F",X"E470",X"F12F",X"008C",X"11B8",X"2059",X"2A4F",X"3041",X"316B",X"2CE9",X"21D1",X"1207",X"00A8",X"F105",X"E3C2",X"D95F",X"D31B",X"D168",X"D4CF",X"DC40",X"E5F2",X"F306",X"03A9",X"14FE",X"2265",X"2BC3",X"314E",X"30EB",X"2ABD",X"1EE4",X"0E4F",X"FCDE",X"EE25",X"E1BF",X"D7B2",X"D26C",X"D207",X"D624",X"DE3C",X"E910",X"F63E",X"0702",X"183A",X"24CE",X"2CC6",X"30D3",X"2F6D",X"27B9",X"1B11",X"0A52",X"F964",X"EB6E",X"E030",X"D758",X"D2B0",X"D35C",X"D8D4",X"E193",X"EC97",X"FA58",X"0B1A",X"1B30",X"2672",X"2D6B",X"2FE8",X"2CC5",X"2414",X"16AC",X"05F2",X"F5E2",X"E8D4",X"DE36",X"D692",X"D372",X"D548",X"DB45",X"E4BB",X"F080",X"FE92",X"0F3C",X"1E00",X"27DD",X"2DCF",X"2F15",X"2AAC",X"20EC",X"12C7",X"01FF",X"F2A0",X"E63C",X"DCB2",X"D671",X"D469",X"D74B",X"DE31",X"E7A5",X"F388",X"024C",X"12B9",X"203B",X"2950",X"2E88",X"2E04",X"2838",X"1D8C",X"0E4F",X"FD8B",X"EF26",X"E3B9",X"DA84",X"D585",X"D54F",X"D8ED",X"E025",X"EA5C",X"F718",X"06C2",X"16A6",X"22BE",X"2AFF",X"2F42",X"2D78",X"2589",X"192A",X"095A",X"F9B2",X"EC7E",X"E192",X"D92F",X"D575",X"D698",X"DB63",X"E321",X"ED9F",X"FAF0",X"0B8A",X"1B0C",X"25C1",X"2C72",X"2F1E",X"2C00",X"22CC",X"14D1",X"0406",X"F4D0",X"E89F",X"DE81",X"D718",X"D45B",X"D6A7",X"DD27",X"E617",X"F0F8",X"FF16",X"0FFA",X"1E8E",X"2809",X"2D96",X"2E4D",X"29A0",X"1F34",X"0FF1",X"FF1A",X"F065",X"E4AA",X"DB61",X"D59A",X"D43A",X"D790",X"DEFA",X"E8C6",X"F48E",X"038D",X"1449",X"217D",X"2A30",X"2EDB",X"2DCB",X"2731",X"1BC8",X"0B97",X"FA8E",X"ECAB",X"E1AA",X"D913",X"D4AA",X"D4F7",X"D96D",X"E1C9",X"ECB2",X"F980",X"08F9",X"18BF",X"24EB",X"2C9F",X"2FBE",X"2D1A",X"24F4",X"17E8",X"0701",X"F678",X"E909",X"DEF4",X"D779",X"D454",X"D61F",X"DC0A",X"E556",X"F0D0",X"FE20",X"0E42",X"1D37",X"27A3",X"2DC0",X"2F42",X"2AE4",X"2102",X"12A0",X"0180",X"F1C4",X"E569",X"DBE8",X"D5D8",X"D45E",X"D7AE",X"DECD",X"E8CD",X"F4C6",X"0320",X"138C",X"20CC",X"2944",X"2E2F",X"2DCC",X"27C7",X"1CB6",X"0D12",X"FC20",X"EDC2",X"E289",X"D9E7",X"D57B",X"D571",X"D9F0",X"E266",X"ED2B",X"F924",X"07CA",X"17A1",X"2378",X"2AB4",X"2DE6",X"2B86",X"240A",X"181A",X"07A1",X"F728",X"EA1D",X"DFE2",X"D840",X"D519",X"D660",X"DC38",X"E5C4",X"F0A4",X"FD33",X"0CAB",X"1B62",X"257D",X"2BB2",X"2DED",X"29F6",X"20F6",X"1430",X"03A6",X"F3CE",X"E77F",X"DE2A",X"D7A3",X"D5B6",X"D87D",X"DF38",X"E8FB",X"F48D",X"01A1",X"10A7",X"1E6F",X"279C",X"2CA6",X"2CDA",X"278D",X"1DE1",X"1015",X"FF60",X"F05F",X"E535",X"DC82",X"D6FC",X"D62E",X"D9CA",X"E147",X"EBC4",X"F75A",X"0456",X"1396",X"20C1",X"2885",X"2C17",X"2B2B",X"2507",X"19E0",X"0AEA",X"FA84",X"EC94",X"E219",X"DA4A",X"D65C",X"D681",X"DAF8",X"E324",X"EDCB",X"F9A7",X"079B",X"1679",X"21D7",X"28BE",X"2B90",X"2912",X"21CE",X"1646",X"06D9",X"F714",X"EA75",X"E0CA",X"D9CC",X"D72E",X"D89B",X"DDE0",X"E6B6",X"F18B",X"FDAC",X"0BC9",X"1976",X"2355",X"299D",X"2B77",X"27A7",X"1F90",X"1370",X"03ED",X"F50A",X"E998",X"E0B2",X"DAC9",X"D94A",X"DB6D",X"E11D",X"E9C4",X"F3F5",X"FFAC",X"0DBF",X"1AA1",X"233D",X"286C",X"2977",X"250E",X"1C82",X"1024",X"00D2",X"F2F6",X"E89F",X"E06E",X"DB37",X"DA77",X"DD0D",X"E2F9",X"EBAB",X"F5B0",X"010D",X"0EAE",X"1AD9",X"22E2",X"277B",X"27F8",X"2300",X"19C0",X"0DA9",X"FED3",X"F1B2",X"E84E",X"E0ED",X"DC8B",X"DBF7",X"DEFA",X"E4ED",X"EDB0",X"F7A1",X"02AB",X"0FC5",X"1B70",X"22C1",X"266F",X"261D",X"20BA",X"1791",X"0B71",X"FD76",X"F124",X"E81B",X"E137",X"DD6C",X"DD85",X"E10D",X"E725",X"EF75",X"F966",X"046C",X"10F3",X"1BFC",X"22D1",X"2604",X"2559",X"1FF1",X"1689",X"0A74",X"FCD8",X"F0E4",X"E811",X"E1A7",X"DE50",X"DE6F",X"E201",X"E83C",X"F054",X"FA01",X"04E1",X"10FA",X"1B2C",X"2182",X"247A",X"239D",X"1E52",X"154E",X"097D",X"FC10",X"EFFC",X"E6AA",X"DFDA",X"DC8B",X"DCC9",X"E028",X"E68E",X"EF15",X"F920",X"044C",X"1124",X"1C2E",X"231E",X"26A8",X"25EC",X"201E",X"168E",X"0A59",X"FC62",X"F02A",X"E6C4",X"E000",X"DCC6",X"DD51",X"E0C7",X"E6C4",X"EEE3",X"F8A2",X"03BF",X"1015",X"1AE7",X"21F0",X"259A",X"2561",X"2048",X"1754",X"0B69",X"FDDE",X"F1DD",X"E88D",X"E193",X"DDF2",X"DDF9",X"E100",X"E692",X"EE5E",X"F7CE",X"01F1",X"0DA1",X"187F",X"1FB6",X"23BA",X"23ED",X"1F9D",X"1758",X"0C75",X"FF9C",X"F382",X"EA14",X"E32A",X"DF6B",X"DF44",X"E1FA",X"E709",X"EE34",X"F706",X"0104",X"0BCA",X"160A",X"1DB3",X"2217",X"22E6",X"1F79",X"1840",X"0E5B",X"02B5",X"F717",X"ED85",X"E684",X"E270",X"E1A3",X"E376",X"E75F",X"ED41",X"F52C",X"FE98",X"08A5",X"1325",X"1BBE",X"212D",X"2330",X"20B7",X"1A62",X"1140",X"05C3",X"F9CD",X"EF5E",X"E773",X"E292",X"E0D9",X"E1EF",X"E528",X"EAC3",X"F261",X"FB5C",X"04E6",X"0F0D",X"180D",X"1E2B",X"213A",X"204D",X"1B47",X"1360",X"0970",X"FE8D",X"F40A",X"EB80",X"E5C7",X"E360",X"E3B2",X"E5B1",X"E9C1",X"EFE3",X"F829",X"0129",X"0A89",X"13AC",X"1ACD",X"1F28",X"1FBE",X"1C5D",X"1614",X"0D93",X"039C",X"F93A",X"F017",X"E96F",X"E5C0",X"E4BF",X"E56B",X"E834",X"ED34",X"F45A",X"FCBE",X"054F",X"0E0A",X"1649",X"1C00",X"1E34",X"1CB2",X"1827",X"114D",X"08AF",X"FED3",X"F514",X"ED54",X"E894",X"E65D",X"E5C6",X"E727",X"EAD9",X"F09F",X"F821",X"0060",X"08A1",X"10C5",X"17B2",X"1BE0",X"1D07",X"1AD8",X"1577",X"0DBD",X"0431",X"FA2A",X"F0CD",X"E979",X"E4F2",X"E2E5",X"E336",X"E5DE",X"EB05",X"F253",X"FAC4",X"038E",X"0CA3",X"1531",X"1B79",X"1E67",X"1DE1",X"19D9",X"12DE",X"0A3D",X"0037",X"F60F",X"EDCC",X"E815",X"E4FD",X"E457",X"E5BB",X"E974",X"EF59",X"F6F2",X"FF62",X"080F",X"104C",X"1719",X"1BF0",X"1DFA",X"1C2A",X"1722",X"0FCF",X"071F",X"FDB2",X"F4A8",X"ED4C",X"E850",X"E632",X"E68C",X"E8C5",X"ED02",X"F31D",X"FA53",X"01E2",X"098B",X"10B0",X"169C",X"1A1C",X"1A66",X"179C",X"123B",X"0B2A",X"02FE",X"FAAF",X"F2DE",X"ED04",X"E984",X"E8ED",X"EA64",X"ED03",X"F108",X"F6AB",X"FD3E",X"03E4",X"0A56",X"1020",X"1426",X"1617",X"1532",X"1167",X"0BB7",X"052A",X"FE43",X"F79B",X"F1F7",X"EEA0",X"EDEF",X"EEFD",X"F109",X"F432",X"F832",X"FD3D",X"02BB",X"07B1",X"0C41",X"1033",X"1279",X"124C",X"1022",X"0C35",X"0706",X"015A",X"FBD6",X"F697",X"F2B1",X"F140",X"F1C7",X"F32D",X"F572",X"F86E",X"FC1D",X"002C",X"0466",X"082B",X"0B8E",X"0DF4",X"0F00",X"0E39",X"0BD8",X"081D",X"036A",X"FE9D",X"F9E4",X"F5CF",X"F313",X"F236",X"F35C",X"F516",X"F709",X"F998",X"FD18",X"00FC",X"04C3",X"0814",X"0A9C",X"0C42",X"0C5B",X"0B1F",X"0844",X"0469",X"005F",X"FCA6",X"F907",X"F5D8",X"F45C",X"F46A",X"F5AA",X"F743",X"F9A7",X"FC5F",X"FF57",X"02CF",X"05F2",X"0851",X"0A12",X"0A9F",X"0A35",X"08B4",X"05F3",X"025B",X"FED7",X"FB82",X"F889",X"F67A",X"F5E9",X"F6B0",X"F819",X"F9F7",X"FC06",X"FE69",X"0142",X"0416",X"05F5",X"07BB",X"0918",X"0955",X"0829",X"05F9",X"033A",X"0022",X"FD23",X"FA0F",X"F7AA",X"F6A2",X"F6CD",X"F814",X"F9DA",X"FB91",X"FD51",X"FF6F",X"01FB",X"0446",X"05F7",X"0757",X"07FB",X"079A",X"0647",X"040D",X"0142",X"FE7C",X"FC24",X"FA33",X"F8ED",X"F87D",X"F922",X"FA72",X"FBB7",X"FD2F",X"FF39",X"016C",X"0363",X"0518",X"065B",X"072F",X"0747",X"0693",X"0509",X"0295",X"003C",X"FE1F",X"FC33",X"FA86",X"F94D",X"F919",X"F9D6",X"FB1A",X"FC6A",X"FDFA",X"FFD0",X"01C3",X"039D",X"04C8",X"0568",X"05E3",X"05BD",X"04DD",X"0341",X"0168",X"FF75",X"FD67",X"FBC8",X"FAA1",X"FA4D",X"FAE0",X"FBDF",X"FCEB",X"FE24",X"FF4F",X"009B",X"0204",X"0386",X"04BB",X"05AC",X"05CB",X"054F",X"045E",X"02CD",X"00FC",X"FF0A",X"FD7F",X"FC66",X"FB9B",X"FB89",X"FC2E",X"FD1B",X"FDEB",X"FE9E",X"FFB5",X"0111",X"0275",X"036B",X"0428",X"04B9",X"04B2",X"0401",X"02BA",X"0162",X"0022",X"FF18",X"FDCC",X"FCC5",X"FC40",X"FC0F",X"FC38",X"FCBF",X"FDBC",X"FEE3",X"0014",X"014F",X"0264",X"031B",X"0378",X"0397",X"0374",X"02A6",X"01A4",X"0067",X"FF58",X"FE22",X"FCF7",X"FC3C",X"FBC9",X"FBD7",X"FC61",X"FD37",X"FE06",X"FEC3",X"FFB3",X"00B9",X"014C",X"01CE",X"0202",X"021C",X"021F",X"01C1",X"00EF",X"FF91",X"FE6F",X"FDDD",X"FD7C",X"FD3B",X"FD25",X"FD6D",X"FE0F",X"FE7E",X"FF4E",X"0004",X"00E8",X"0192",X"0208",X"025E",X"0294",X"02A4",X"0237",X"0164",X"007D",X"FF99",X"FEE9",X"FE70",X"FE1B",X"FE3F",X"FE91",X"FED3",X"FF11",X"FF89",X"0021",X"00C6",X"0124",X"0177",X"01D7",X"020B",X"0202",X"01C7",X"011C",X"0057",X"FFC4",X"FF2A",X"FE98",X"FE48",X"FE1A",X"FE1B",X"FE36",X"FE67",X"FEE2",X"FF79",X"002D",X"0091",X"00E4",X"0120",X"012D",X"0141",X"012C",X"00A3",X"0035",X"FFD4",X"FF61",X"FEDB",X"FE7E",X"FE9A",X"FEE4",X"FF28",X"FFA2",X"0002",X"0027",X"004E",X"00D4",X"0132",X"0197",X"01E3",X"01E6",X"01C7",X"016D",X"00DC",X"0022",X"FFA8",X"FF46",X"FF03",X"FEDA",X"FF06",X"FF34",X"FF70",X"FFDD",X"FFFA",X"FFF3",X"0035",X"00B3",X"0168",X"01A8",X"0172",X"0134",X"00BC",X"0017",X"FFAB",X"FF1C",X"FEEE",X"FF1E",X"FF81",X"FFA0",X"FFBF",X"FFE5",X"FFFD",X"0023",X"0094",X"0108",X"0161",X"0180",X"0174",X"0177",X"014C",X"00F5",X"0084",X"0028",X"FFC6",X"FF5A",X"FF33",X"FF1C",X"FEFA",X"FEFB",X"FF28",X"FF8C",X"FFCB",X"000E",X"005B",X"0087",X"00A3",X"0093",X"008B",X"0099",X"006C",X"002E",X"FFE8",X"FF49",X"FEC6",X"FE8E",X"FE3E",X"FE0C",X"FE29",X"FE76",X"FEDD",X"FF33",X"FF8B",X"FFF3",X"001E",X"003D",X"006D",X"0099",X"00AB",X"00C4",X"00A3",X"003F",X"FFCE",X"FF70",X"FF24",X"FEE0",X"FEBB",X"FED5",X"FEC5",X"FEFD",X"FF52",X"FF93",X"FFB0",X"FFEE",X"0055",X"006E",X"0093",X"00AC",X"0098",X"0034",X"FFE9",X"FF61",X"FEDF",X"FE62",X"FE4F",X"FE63",X"FEAA",X"FEBE",X"FEED",X"FF2D",X"FF8C",X"FFEF",X"0040",X"00C5",X"010D",X"0118",X"0147",X"00FC",X"009F",X"0083",X"002A",X"FFB6",X"FF89",X"FF46",X"FF23",X"FF0E",X"FF46",X"FF95",X"FFDA",X"0008",X"0040",X"007D",X"00C2",X"0100",X"015D",X"0171",X"0161",X"00FA",X"0094",X"0025",X"FFA3",X"FF71",X"FF83",X"FF3B",X"FF3D",X"FF19",X"FF17",X"FF58",X"FFBF",X"0030",X"007C",X"00DB",X"011C",X"0193",X"01AE",X"017A",X"012C",X"00BC",X"003F",X"0000",X"FFB9",X"FF37",X"FEE1",X"FE86",X"FE88",X"FE9B",X"FEED",X"FF6D",X"FFEE",X"005B",X"00E3",X"0132",X"0177",X"01C1",X"0198",X"0175",X"0166",X"00D3",X"0064",X"0012",X"FFAA",X"FF92",X"FF2B",X"FF1E",X"FEEA",X"FF2D",X"FFB1",X"001B",X"00B4",X"0107",X"0129",X"0174",X"016A",X"0139",X"00EE",X"00C9",X"0082",X"001F",X"FFC8",X"FF4C",X"FED1",X"FE6A",X"FE80",X"FE82",X"FECF",X"FEC5",X"FF1A",X"FF9C",X"001B",X"0039",X"0055",X"0099",X"00C6",X"00AB",X"0082",X"0039",X"FFD7",X"FF9F",X"FF98",X"FF42",X"FF1B",X"FED7",X"FED6",X"FEE7",X"FEF4",X"FF3F",X"FFA0",X"FFE2",X"0016",X"0070",X"00C7",X"00E0",X"011B",X"0111",X"00D7",X"009A",X"0065",X"001D",X"FFAF",X"FF54",X"FF1F",X"FEF9",X"FEED",X"FED9",X"FEEA",X"FF2B",X"FFCB",X"0016",X"0040",X"0051",X"004C",X"003C",X"006D",X"009B",X"00AC",X"0064",X"0005",X"FF75",X"FF2C",X"FF25",X"FEFB",X"FEB0",X"FE87",X"FED8",X"FF13",X"FF33",X"FF9E",X"FFE3",X"0011",X"003A",X"0097",X"0084",X"007F",X"0095",X"008F",X"003A",X"FFBF",X"FF74",X"FF28",X"FEFE",X"FF13",X"FF4F",X"FF7A",X"FF9D",X"FFBD",X"FFFD",X"0000",X"000F",X"003E",X"0090",X"00B5",X"00AE",X"0099",X"007A",X"004D",X"0027",X"001F",X"000D",X"FFC3",X"FFCA",X"FFE2",X"FFF5",X"FFEC",X"000F",X"0024",X"0048",X"0073",X"00BE",X"011C",X"012A",X"013F",X"0172",X"0154",X"0118",X"00D0",X"009E",X"0087",X"003E",X"001C",X"0021",X"002F",X"000B",X"FFF9",X"FFFA",X"FFFF",X"0016",X"0055",X"0057",X"0041",X"0062",X"0073",X"0071",X"0067",X"0032",X"FFF6",X"FFD1",X"FFBA",X"FFA8",X"FF8D",X"FF5F",X"FF7F",X"FF87",X"FF76",X"FF8C",X"FF9D",X"FFA2",X"FFCC",X"FFCB",X"FFA2",X"FF87",X"FF97",X"FF7C",X"FF62",X"FF21",X"FF11",X"FF06",X"FF32",X"FF3C",X"FF57",X"FF4B",X"FF88",X"FFB3",X"FFE3",X"0014",X"005D",X"0086",X"00C0",X"00D8",X"00E2",X"00AA",X"0097",X"0097",X"009A",X"0083",X"004D",X"FFF0",X"FFD7",X"FFFE",X"FFED",X"FFB8",X"FFA4",X"FF94",X"FF90",X"FFBA",X"FFCC",X"FFE9",X"FFF7",X"0000",X"FFC5",X"FFAD",X"FFC7",X"FFC6",X"FFA6",X"FF93",X"FFA6",X"FF9F",X"FF71",X"FF5B",X"FF45",X"FF5A",X"FF8B",X"FFD7",X"0001",X"001A",X"0040",X"0047",X"0033",X"002F",X"004D",X"001D",X"000C",X"FFFF",X"FFC4",X"FF9C",X"FF80",X"FF6B",X"FF45",X"FF45",X"FF72",X"FFA6",X"FFA7",X"FF81",X"FF76",X"FF47",X"FF48",X"FF7F",X"FF98",X"FFEF",X"003C",X"0024",X"FFEA",X"FFCC",X"FFD6",X"FFD0",X"FFBA",X"FFC0",X"FFF8",X"0013",X"0009",X"FFED",X"FFDA",X"FFEE",X"000E",X"002E",X"005F",X"0092",X"00A0",X"00B1",X"0096",X"0088",X"0083",X"007E",X"0071",X"005D",X"007D",X"00AD",X"0095",X"00A7",X"00B1",X"008B",X"0087",X"008E",X"00F3",X"011D",X"011C",X"011A",X"00DC",X"00A8",X"008A",X"004C",X"0052",X"0084",X"0096",X"00AC",X"0067",X"0050",X"000D",X"FFE2",X"FFCC",X"FFBA",X"FFC6",X"FFC8",X"FFB4",X"FFC3",X"FFBE",X"FFAF",X"FFEF",X"0017",X"FFF7",X"FFEE",X"FFF7",X"FFFE",X"0018",X"FFFD",X"FFBF",X"FFA4",X"FFB6",X"FFBD",X"FFD8",X"FFD1",X"FFA4",X"FF77",X"FF75",X"FF84",X"FF93",X"FFB2",X"FFCE",X"FFEB",X"FFC8",X"FFB4",X"FFD8",X"FFC0",X"FFDB",X"FFD5",X"FFE2",X"FFA1",X"FF7B",X"FF68",X"FF8C",X"FF88",X"FF9D",X"FF82",X"FFBB",X"0001",X"0017",X"FFFB",X"FFF5",X"000A",X"FFF9",X"FFBF",X"FF8D",X"FF87",X"FFA7",X"FFAD",X"FF9C",X"FF95",X"FFB2",X"FFBA",X"FFFD",X"0017",X"000E",X"FFED",X"FFFA",X"0009",X"0023",X"0046",X"0056",X"0070",X"006A",X"0060",X"004D",X"0044",X"005A",X"005E",X"002A",X"0010",X"FFFF",X"FFC3",X"FF72",X"FF44",X"FF56",X"FF4E",X"FF50",X"FF6E",X"FF80",X"FF86",X"FF7C",X"FF7F",X"FFAB",X"FFBA",X"FFD8",X"FFA6",X"FFA9",X"FFCA",X"FFEF",X"FFB4",X"FF85",X"FF55",X"FF33",X"FF5A",X"FFA6",X"FFAA",X"FF7E",X"FF78",X"FF8E",X"FFB2",X"FFC2",X"FFD7",X"FFFC",X"0044",X"006F",X"0069",X"004C",X"004D",X"0036",X"005D",X"0091",X"0077",X"0060",X"004A",X"0052",X"0072",X"003D",X"0014",X"0023",X"0038",X"0071",X"006B",X"002B",X"0035",X"0044",X"0047",X"0068",X"0085",X"008B",X"0085",X"0095",X"0099",X"007D",X"0078",X"0076",X"0057",X"0020",X"0000",X"0019",X"0004",X"000C",X"003D",X"0040",X"0032",X"001A",X"FFF0",X"FFAC",X"FF94",X"FFC3",X"FFF6",X"FFE1",X"FFE0",X"FFE0",X"FFEB",X"FFF6",X"FFFD",X"0020",X"0007",X"0037",X"001A",X"0019",X"0008",X"001E",X"0027",X"0018",X"002D",X"0002",X"0015",X"002B",X"FFFC",X"FFFF",X"FFF7",X"FFB3",X"FF80",X"FF55",X"FF6D",X"FFB1",X"FFCA",X"FFC7",X"FFA5",X"FF64",X"FF63",X"FF86",X"FF9C",X"FFD5",X"0004",X"0007",X"FFF2",X"FFE6",X"FFE7",X"FFC2",X"FFC6",X"FFEA",X"0007",X"FFEF",X"FFD8",X"FFCF",X"FFDA",X"FFCA",X"FFBF",X"FFD8",X"FFDB",X"FFCB",X"FFD3",X"FFC3",X"FFBE",X"FFB7",X"FFA9",X"FF82",X"FF3D",X"FF31",X"FF55",X"FF81",X"FFB4",X"FFF5",X"0009",X"FFB5",X"FF78",X"FF74",X"FF9D",X"FFBB",X"FFD7",X"FFC7",X"FFC6",X"0000",X"0005",X"FFEF",X"FFBD",X"FFC7",X"FFDF",X"0012",X"0021",X"001F",X"FFFA",X"FFFF",X"FFFC",X"FFE3",X"FFDA",X"000A",X"0019",X"000B",X"FFF3",X"0003",X"FFF4",X"FFD9",X"FFEB",X"FFFB",X"FFF1",X"0004",X"0027",X"0048",X"0058",X"005A",X"0068",X"005A",X"0068",X"0098",X"00C7",X"00C8",X"00BA",X"00AA",X"00A3",X"006A",X"007F",X"007B",X"0084",X"0084",X"0051",X"0043",X"0022",X"000D",X"FFE2",X"FFCB",X"FFD4",X"FFEF",X"FFED",X"FFB7",X"FF99",X"FFAF",X"000E",X"0047",X"003F",X"007B",X"00C1",X"009F",X"0080",X"0058",X"001B",X"001E",X"001D",X"0017",X"002C",X"0015",X"FFE9",X"FFB7",X"FFB0",X"FF98",X"FFC7",X"FFF8",X"FFF0",X"0006",X"001B",X"002D",X"0056",X"0050",X"004A",X"004C",X"0067",X"004E",X"0028",X"0014",X"FFF1",X"FFCC",X"FFB8",X"FFDB",X"FFF0",X"0006",X"0011",X"0001",X"0014",X"0043",X"0036",X"0022",X"0020",X"0028",X"002F",X"0009",X"FFEB",X"FFB0",X"FFAA",X"FFBF",X"FFAD",X"FF7C",X"FF63",X"FF5B",X"FF5C",X"FF1D",X"FF25",X"FF2C",X"FF34",X"FF3A",X"FF46",X"FF72",X"FF83",X"FF97",X"FFB4",X"FFE4",X"FFD8",X"FFD2",X"FFDA",X"FFA2",X"FF82",X"FFB0",X"FFD6",X"FFFE",X"FFEC",X"FFC4",X"FFC3",X"FFD0",X"FFD4",X"FFB0",X"FF95",X"FFA6",X"FFAB",X"FFAD",X"FFAB",X"FF99",X"FF4A",X"FF25",X"FF26",X"FF2E",X"FF36",X"FF3E",X"FF6D",X"FF89",X"FF9C",X"FFAF",X"FFD5",X"FFA1",X"FF95",X"FFD3",X"0006",X"0013",X"FFF7",X"FFF3",X"FFF2",X"FFE7",X"FFFA",X"0001",X"0010",X"FFF1",X"FFE6",X"FFFD",X"FFE7",X"0000",X"0024",X"001A",X"003C",X"0077",X"00A9",X"007C",X"005B",X"0072",X"006A",X"0094",X"0097",X"005D",X"0021",X"FFF5",X"FFF5",X"0004",X"0012",X"0013",X"001B",X"0008",X"001F",X"003C",X"0059",X"0075",X"009A",X"008A",X"009D",X"00C2",X"00D0",X"00A4",X"0062",X"003D",X"0008",X"0008",X"005A",X"0070",X"0085",X"0088",X"0089",X"005E",X"0030",X"002C",X"0061",X"0090",X"006B",X"0003",X"FF99",X"FFB6",X"FFC7",X"FFCD",X"FFC4",X"FFE6",X"FFC6",X"FFA1",X"FF84",X"FF92",X"FFAE",X"FFAC",X"FF86",X"FF8B",X"FF86",X"FFA7",X"FF96",X"FFAE",X"FFB8",X"FF99",X"FF6C",X"FF68",X"FF62",X"FF88",X"FFA6",X"FF9C",X"FF7B",X"FF72",X"FF90",X"FFF7",X"0019",X"001B",X"0029",X"0034",X"0039",X"0054",X"0087",X"00BF",X"00EC",X"00E5",X"00CC",X"00B4",X"00A5",X"008B",X"00A2",X"00C4",X"00F9",X"00B9",X"0080",X"0076",X"005E",X"005A",X"0020",X"0000",X"FFFE",X"000E",X"0011",X"0022",X"0050",X"0037",X"FFF2",X"FFA3",X"FF95",X"FF9E",X"FF90",X"FF4F",X"FF33",X"FF34",X"FF36",X"FF14",X"FF11",X"FF23",X"FF30",X"FF61",X"FF82",X"FF71",X"FF5D",X"FF4B",X"FF35",X"FF21",X"FF45",X"FF32",X"FF18",X"FEEC",X"FEEC",X"FEE3",X"FEEF",X"FEF7",X"FF05",X"FF22",X"FF6D",X"FFC1",X"FFFD",X"FFED",X"FFED",X"0025",X"002F",X"0019",X"0048",X"0057",X"0070",X"0060",X"0052",X"0065",X"006A",X"0052",X"0064",X"0089",X"009B",X"00AD",X"00B0",X"00B4",X"0085",X"0039",X"007D",X"00C8",X"00AA",X"007B",X"004F",X"0074",X"008B",X"0087",X"0091",X"00BA",X"00BD",X"009B",X"0094",X"0099",X"0091",X"0093",X"0087",X"00AA",X"00AA",X"00A3",X"00B2",X"0099",X"007C",X"006C",X"003C",X"0013",X"FFF9",X"FFE6",X"FFDB",X"FFEF",X"FFD9",X"FFAD",X"FF7D",X"FF44",X"FF19",X"FEF9",X"FF39",X"FF6A",X"FF5E",X"FF5D",X"FF60",X"FF78",X"FF9D",X"FF94",X"FF82",X"FF5A",X"FF65",X"FF7E",X"FF9B",X"FF9D",X"FFAB",X"FFB7",X"FFB0",X"FFBA",X"FFDD",X"0005",X"0035",X"0069",X"006A",X"0090",X"009D",X"0076",X"0048",X"004E",X"0061",X"0083",X"0076",X"0070",X"005B",X"0061",X"0060",X"0050",X"0049",X"0043",X"0040",X"0020",X"0001",X"FFF2",X"FFE6",X"FFD0",X"FF9D",X"FF58",X"FF40",X"FF30",X"FF6E",X"FF71",X"FF60",X"FF5E",X"FF58",X"FF31",X"FF24",X"FF3E",X"FF6D",X"FF8F",X"FFCC",X"000E",X"0022",X"0003",X"FFFE",X"002C",X"0026",X"FFFC",X"FFDD",X"FFD9",X"FFD4",X"FFD5",X"FFDA",X"FFDF",X"FF73",X"FF5A",X"FF8D",X"FFB9",X"FFC5",X"FFDA",X"FFCB",X"FFD0",X"FFBB",X"FF5E",X"FF79",X"FFA1",X"FFFB",X"001C",X"000D",X"FFF2",X"FFB7",X"FF9E",X"FFBE",X"FFDA",X"FFEC",X"FFE0",X"FFE5",X"0007",X"FFE3",X"FFED",X"FFEE",X"FFEC",X"FFE3",X"FFFC",X"FFFA",X"0005",X"0005",X"000B",X"002E",X"0017",X"FFFD",X"0010",X"0016",X"FFFB",X"FFDD",X"FFFB",X"FFF9",X"FFFE",X"FFFE",X"000F",X"0015",X"0028",X"0069",X"0065",X"0054",X"0065",X"0060",X"0051",X"007F",X"0097",X"00A1",X"0083",X"006A",X"007D",X"009E",X"00AF",X"00BD",X"00B1",X"00BC",X"00A1",X"009D",X"0079",X"0036",X"0034",X"0031",X"0002",X"FFE6",X"FFC8",X"FFB9",X"FFA7",X"FFA3",X"FF87",X"FFA1",X"FFD4",X"0000",X"0003",X"0007",X"0036",X"0016",X"0006",X"001B",X"0047",X"0042",X"003F",X"0043",X"001D",X"0006",X"FFDE",X"FFBB",X"FF9F",X"FFB9",X"FFE4",X"0032",X"0032",X"0024",X"000A",X"000B",X"000F",X"0025",X"004D",X"0032",X"0052",X"007E",X"0093",X"0091",X"0049",X"0043",X"0031",X"FFFE",X"0003",X"FFF3",X"FFDF",X"FFDA",X"FFB7",X"FF94",X"FF6E",X"FF58",X"FF74",X"FF85",X"FFA0",X"FFB9",X"FFDE",X"FFD3",X"FFC7",X"FFC7",X"FFCA",X"FFBE",X"FF97",X"FF90",X"FFBE",X"FFF6",X"FFE1",X"FFCC",X"FF9B",X"FF7F",X"FF7E",X"FF8A",X"FF8B",X"FFAD",X"FFBC",X"FFAD",X"FFA5",X"FF89",X"FF6C",X"FF54",X"FF49",X"FF6F",X"FF83",X"FF95",X"FF85",X"FF52",X"FF51",X"FF68",X"FF63",X"FF6C",X"FF84",X"FFB8",X"FFE8",X"0005",X"FFDE",X"FF94",X"FF98",X"FFD9",X"0001",X"FFF5",X"0005",X"0005",X"FFFE",X"FFF1",X"FFE5",X"FFE5",X"000C",X"004C",X"0086",X"00A9",X"00A0",X"0074",X"0062",X"0083",X"007D",X"006C",X"0056",X"004D",X"0075",X"005C",X"000C",X"FFF3",X"FFE7",X"FFF0",X"001F",X"0028",X"0029",X"0064",X"0027",X"FFDE",X"FFF0",X"0020",X"0070",X"0072",X"0055",X"0031",X"FFEC",X"FFF1",X"FFED",X"FFDE",X"FFC4",X"FFCB",X"FFA3",X"FF84",X"FF92",X"FF8F",X"FF8D",X"FFAE",X"FF9C",X"FFB2",X"FFC0",X"FFDC",X"FFDB",X"FFFA",X"0003",X"FFE5",X"FFFE",X"0016",X"001A",X"006C",X"0091",X"007A",X"006F",X"005E",X"0061",X"0085",X"0082",X"005E",X"004E",X"0053",X"0059",X"003E",X"003B",X"0050",X"0062",X"0050",X"0031",X"0010",X"001A",X"0054",X"0082",X"0095",X"00A8",X"00A5",X"0090",X"009C",X"00A0",X"0061",X"0002",X"FFC4",X"FFBB",X"FFA4",X"FFB0",X"FFDC",X"FFEB",X"FFBB",X"FFB5",X"FF98",X"FFA6",X"FFB5",X"FFB5",X"FFA7",X"FF84",X"FF61",X"FF56",X"FF70",X"FFA1",X"FF98",X"FF81",X"FF54",X"FF45",X"FF94",X"FFA8",X"FF74",X"FF78",X"FFB3",X"FFBE",X"FFA1",X"FFA7",X"FFB1",X"FFB6",X"FF9E",X"FFA6",X"FF8B",X"FF8B",X"FFD1",X"000F",X"0041",X"0026",X"FFD3",X"FF74",X"FF50",X"FF50",X"FF80",X"FFA6",X"FF8B",X"FF87",X"FF94",X"FFB1",X"FF89",X"FF45",X"FF5E",X"FF84",X"FF8F",X"FFC9",X"FFE9",X"0004",X"001E",X"001F",X"0015",X"0022",X"0024",X"0030",X"004D",X"0075",X"008E",X"008B",X"008D",X"0097",X"00B8",X"00A8",X"00C5",X"00D9",X"00CB",X"00C4",X"006F",X"0020",X"FFF5",X"FFF3",X"0038",X"0066",X"0056",X"FFFD",X"FFBE",X"FFB0",X"FFC6",X"FFB5",X"FFB2",X"FFCC",X"000F",X"001B",X"0063",X"007B",X"009D",X"00BE",X"00D0",X"00A2",X"0070",X"0056",X"004A",X"003B",X"0057",X"004D",X"003E",X"0015",X"FFF6",X"FFD7",X"FFB3",X"FFAE",X"FFD4",X"FFF5",X"FFFD",X"0002",X"000F",X"0020",X"0000",X"000D",X"FFF9",X"FFF5",X"FFE5",X"FFF6",X"FFF8",X"FFA7",X"FF56",X"FF41",X"FF6A",X"FF87",X"FFAE",X"FFD5",X"FFE1",X"FFBB",X"FF9E",X"FF9D",X"FFB9",X"FFC7",X"FFE0",X"0019",X"003F",X"0045",X"0010",X"FFF7",X"0003",X"0029",X"0030",X"0054",X"008D",X"0096",X"00A8",X"0091",X"003B",X"001E",X"0026",X"000B",X"0009",X"0054",X"0085",X"00A8",X"0089",X"0043",X"0038",X"0037",X"0045",X"0029",X"0017",X"0022",X"0020",X"FFE8",X"FFC8",X"FFCD",X"FFB4",X"FF99",X"FF56",X"FF2E",X"FF2D",X"FF3D",X"FF53",X"FF57",X"FF58",X"FF45",X"FF44",X"FF19",X"FF14",X"FF48",X"FF99",X"FFC2",X"FFA4",X"FF86",X"FF75",X"FF82",X"FFA7",X"FF99",X"FF8E",X"FF78",X"FF92",X"FFA2",X"FFB1",X"FF7A",X"FF5E",X"FF58",X"FF23",X"FF38",X"FF8A",X"FF96",X"FF9D",X"FF92",X"FF63",X"FF84",X"FFCD",X"0009",X"0021",X"0028",X"002D",X"000E",X"FFFA",X"FFF7",X"FFF9",X"FFF3",X"001A",X"002D",X"001F",X"0000",X"FFED",X"FFFF",X"0008",X"0002",X"0011",X"001A",X"0009",X"000E",X"004D",X"0067",X"0046",X"0045",X"0015",X"0028",X"0056",X"004A",X"0069",X"0079",X"0070",X"0030",X"0020",X"0056",X"0066",X"003A",X"003D",X"0071",X"0074",X"0038",X"000B",X"FFF0",X"FFFD",X"FFFA",X"001A",X"0045",X"0042",X"0074",X"0067",X"0067",X"005D",X"0062",X"002F",X"FFEC",X"FFE0",X"0000",X"0028",X"FFF4",X"FFD4",X"FFA6",X"FF7D",X"FF7B",X"FF8B",X"FF8D",X"FF6E",X"FF6F",X"FFB1",X"FFE4",X"FFF2",X"FFF7",X"000C",X"0046",X"005C",X"007F",X"008B",X"00AD",X"00C1",X"00C2",X"006F",X"0061",X"009C",X"00D5",X"00AB",X"0079",X"003D",X"004B",X"0092",X"0099",X"0072",X"003F",X"0020",X"0039",X"0038",X"000F",X"FFF6",X"FFFE",X"0003",X"FFF1",X"FFDB",X"FFD9",X"FFAE",X"FF8B",X"FF9D",X"FFB8",X"FFA3",X"FF5C",X"FF2C",X"FF25",X"FF37",X"FF49",X"FF24",X"FF41",X"FF6B",X"FF4B",X"FF18",X"FF11",X"FF06",X"FF20",X"FF34",X"FF50",X"FF86",X"FFD8",X"0013",X"0037",X"0037",X"0033",X"0038",X"0018",X"004B",X"0054",X"005A",X"0047",X"0048",X"0028",X"0002",X"FFDC",X"001C",X"0024",X"002A",X"000E",X"000D",X"FFF2",X"FFE0",X"FFEA",X"FFEC",X"FFD0",X"FFDF",X"000F",X"001F",X"0005",X"FFE5",X"FFB2",X"FFA4",X"FFC2",X"FFE3",X"FFD0",X"FFBD",X"FF88",X"FF84",X"FF72",X"FF6F",X"FF6D",X"FF87",X"FFA6",X"FFE2",X"0011",X"0031",X"0038",X"0022",X"001E",X"005C",X"006E",X"0079",X"006C",X"0040",X"0039",X"0039",X"0062",X"004A",X"003A",X"0027",X"0028",X"0047",X"002B",X"002B",X"0006",X"0002",X"0008",X"000C",X"0004",X"002D",X"002A",X"0029",X"0034",X"FFF8",X"FFFA",X"FFD9",X"FFF3",X"FFFF",X"001A",X"0025",X"0008",X"FFDC",X"000B",X"FFF6",X"FFE0",X"FFE8",X"FFF9",X"FFDF",X"FFC5",X"FFCA",X"FFDF",X"FFCD",X"FFE2",X"FFEF",X"FFFB",X"FFFB",X"FFEE",X"FFCF",X"FFD1",X"FFE8",X"0016",X"0032",X"0056",X"0048",X"0013",X"FFF7",X"FFFF",X"0027",X"006D",X"007D",X"0052",X"0047",X"0062",X"0087",X"007B",X"0050",X"0043",X"0063",X"0080",X"006C",X"0072",X"0054",X"0039",X"0032",X"0017",X"001B",X"0011",X"0001",X"0002",X"FFE0",X"FFB4",X"FF9C",X"FFAA",X"FFC9",X"FFC2",X"FFD9",X"FFF0",X"FFD1",X"FFA8",X"FFD4",X"FFBA",X"FF88",X"FF84",X"FFA4",X"FFC4",X"FFD2",X"FFCA",X"FFB1",X"FFA0",X"FF92",X"FF62",X"FF7B",X"FFCE",X"FFDD",X"FFC9",X"FF9F",X"FF7D",X"FF68",X"FF46",X"FF2B",X"FF51",X"FF76",X"FF7F",X"FF93",X"FF61",X"FF1B",X"FF22",X"FF28",X"FF4A",X"FF4D",X"FF94",X"FFBD",X"FFA5",X"FF9F",X"FF9A",X"FF97",X"FFB3",X"FFDB",X"FFE8",X"FFF2",X"0005",X"FFFF",X"FFF7",X"FFDD",X"FFE5",X"FFDA",X"FFDC",X"0009",X"0032",X"0066",X"0070",X"005D",X"003A",X"001D",X"0044",X"006B",X"0078",X"006B",X"0038",X"0042",X"003C",X"0040",X"0041",X"0058",X"007C",X"006D",X"0069",X"006B",X"0044",X"000B",X"FFD5",X"000B",X"0018",X"0017",X"0035",X"0012",X"FFD1",X"FFB6",X"FFBB",X"FF9B",X"FFA3",X"FFB1",X"FFE0",X"FFDC",X"FFC7",X"FFB0",X"FFA6",X"FF8B",X"FF70",X"FFB7",X"FFE9",X"000D",X"0008",X"0013",X"0017",X"0047",X"006E",X"009C",X"0066",X"0054",X"008D",X"00C0",X"00E6",X"010A",X"0115",X"00E0",X"0095",X"007C",X"001E",X"FFEE",X"FFED",X"0014",X"000D",X"FFF6",X"0001",X"000B",X"0034",X"0064",X"0085",X"0071",X"0046",X"003A",X"0064",X"008C",X"008B",X"0099",X"007D",X"0063",X"0071",X"0060",X"003D",X"000E",X"FFDF",X"FFE2",X"FFEF",X"FFCE",X"FFCB",X"FFDB",X"FFEC",X"FFE1",X"FFC4",X"FFA0",X"FF93",X"FF90",X"FF7F",X"FF8E",X"FF6D",X"FF61",X"FFA6",X"FFC3",X"FFF6",X"001A",X"FFFF",X"FFBE",X"FFB3",X"FFF2",X"FFE2",X"FFD0",X"FFD6",X"0012",X"001B",X"FFF9",X"FFC7",X"FF9D",X"FF99",X"FF80",X"FF7D",X"FF89",X"FFAE",X"FFA1",X"FFB4",X"FF98",X"FF4C",X"FF2C",X"FF44",X"FF46",X"FF59",X"FF5F",X"FF6B",X"FF89",X"FF86",X"FF8B",X"FF83",X"FF84",X"FFD2",X"0017",X"FFFD",X"FFF4",X"0000",X"FFDD",X"FFE6",X"0015",X"0038",X"0039",X"FFFB",X"FFFF",X"0009",X"000D",X"001B",X"003F",X"0029",X"002F",X"0032",X"FFE6",X"FFC3",X"FFD6",X"FFCF",X"FFD5",X"FFE4",X"FFE8",X"FFE7",X"FFDB",X"FFD7",X"FFDA",X"FFFB",X"0013",X"FFDE",X"FFE4",X"FFCB",X"FFDE",X"FFF5",X"FFFB",X"FFF4",X"FFCE",X"FFAD",X"FFD1",X"FFC1",X"FFEE",X"0012",X"0041",X"004C",X"0053",X"0036",X"0053",X"005E",X"0052",X"0051",X"0041",X"0051",X"005A",X"007B",X"009D",X"0080",X"0061",X"0069",X"0078",X"0032",X"0013",X"000A",X"0023",X"0037",X"0058",X"0017",X"FFA6",X"FF8B",X"FFC9",X"FFD8",X"FFE0",X"FFD9",X"FFFF",X"FFFA",X"000E",X"0013",X"FFEE",X"0001",X"FFF8",X"FFFA",X"FFFE",X"FFD5",X"FFC8",X"FFDC",X"001F",X"0025",X"0030",X"0047",X"005B",X"006C",X"006D",X"0073",X"004F",X"004B",X"0045",X"003D",X"FFFC",X"FFF7",X"FFFE",X"0001",X"FFFF",X"0032",X"0033",X"0002",X"0003",X"0012",X"002D",X"003A",X"000F",X"FFDA",X"FFB4",X"FFB9",X"FFD7",X"FFCF",X"FFBA",X"FF7D",X"FF96",X"FFD4",X"FFE3",X"FFD7",X"FFB6",X"FF96",X"FF73",X"FF74",X"FF4F",X"FF60",X"FFA3",X"FFCA",X"FFBD",X"FF98",X"FFA2",X"FF80",X"FF53",X"FF4B",X"FF64",X"FF73",X"FF71",X"FF69",X"FF53",X"FF4E",X"FF69",X"FF94",X"FF96",X"FF84",X"FF85",X"FF9E",X"FFCF",X"FFEB",X"0009",X"0015",X"001C",X"0034",X"0034",X"0052",X"005F",X"006E",X"0059",X"001A",X"FFEE",X"FFF9",X"000A",X"0009",X"0011",X"0032",X"0021",X"0028",X"003C",X"0047",X"002C",X"0029",X"0025",X"FFF9",X"0011",X"0041",X"003A",X"0012",X"FFEF",X"FFE6",X"FFC0",X"FFBD",X"FFDB",X"FFF3",X"FFF6",X"0001",X"FFE4",X"FFD9",X"FFA2",X"FF8A",X"FFA5",X"FFE2",X"003D",X"0068",X"0049",X"0027",X"0011",X"0007",X"0008",X"003A",X"0041",X"0034",X"0013",X"0009",X"FFC0",X"FFA1",X"FFA2",X"FFA9",X"FFE8",X"003A",X"004E",X"0048",X"0030",X"002A",X"0007",X"FFD9",X"0003",X"003E",X"0076",X"009F",X"00CA",X"00CF",X"00D2",X"0091",X"0045",X"0040",X"006C",X"0091",X"00A8",X"0093",X"008F",X"0072",X"005A",X"0041",X"004A",X"004D",X"0055",X"005C",X"009C",X"009C",X"0071",X"FFF6",X"FFB2",X"FFDD",X"0009",X"0024",X"0015",X"0019",X"001D",X"002B",X"FFFC",X"FFF6",X"FFCF",X"FFC5",X"FFCD",X"FFDC",X"FFD3",X"FFBE",X"FFB2",X"FFA3",X"FFBB",X"FFBC",X"FFE0",X"FFE9",X"FFE7",X"FFEE",X"FFEE",X"FFCA",X"FFA4",X"FF83",X"FF50",X"FF1F",X"FF33",X"FF58",X"FFA8",X"FFBA",X"FF9E",X"FF4E",X"FF3F",X"FF1D",X"FF5C",X"FF55",X"FF34",X"FF4A",X"FF5F",X"FF60",X"FF49",X"FF39",X"FF6B",X"FF97",X"FFA5",X"FFCB",X"FFDA",X"FFCC",X"FFC0",X"FFE7",X"FFDB",X"FFFB",X"002D",X"0075",X"005C",X"0037",X"0027",X"0013",X"0013",X"0011",X"0038",X"0059",X"006C",X"004C",X"002E",X"0015",X"0004",X"0013",X"0004",X"FFFE",X"FFF1",X"000E",X"FFF5",X"FFF2",X"FFEC",X"FFB2",X"FF95",X"FFB6",X"0000",X"FFFE",X"FFD6",X"0000",X"0021",X"FFED",X"FF89",X"FF73",X"FF7B",X"FF9B",X"FFD2",X"FFE3",X"FFB9",X"FFA2",X"FFA8",X"FF96",X"FFBD",X"FF8F",X"FFAA",X"FFCD",X"FFF9",X"FFDA",X"FFCE",X"FFD3",X"000B",X"004B",X"0061",X"0052",X"0035",X"0021",X"003A",X"004F",X"0016",X"001D",X"FFF3",X"0001",X"0013",X"0036",X"0029",X"0030",X"0005",X"0004",X"0011",X"003D",X"0055",X"0059",X"0067",X"0059",X"0065",X"0066",X"0081",X"0065",X"006B",X"007E",X"0080",X"009A",X"0063",X"0041",X"0024",X"001F",X"0043",X"0055",X"0040",X"004F",X"0087",X"0095",X"0079",X"003F",X"0022",X"0031",X"0078",X"004F",X"001E",X"0008",X"0002",X"0001",X"0005",X"FFCF",X"FFD4",X"FFE0",X"FFE1",X"FFBD",X"FFB7",X"FF8F",X"FF77",X"FF6A",X"FF7C",X"FF8A",X"FF80",X"FF7B",X"FF8D",X"FF63",X"FF88",X"FFB8",X"FFC7",X"FFFC",X"FFDF",X"FFC7",X"FFEE",X"0001",X"FFE2",X"FF9F",X"FF97",X"FFBC",X"FFCC",X"FFDD",X"FFF7",X"FFDC",X"FFDE",X"FFFF",X"0001",X"FFE9",X"FFFD",X"FFFF",X"FFF4",X"FFF9",X"000A",X"0044",X"0035",X"0005",X"000E",X"0017",X"0019",X"FFFC",X"FFE7",X"FF9D",X"FFB5",X"FFD7",X"FFFA",X"FFD3",X"FFA6",X"FF88",X"FF85",X"FF98",X"FF8B",X"FF96",X"FFA5",X"FFB5",X"FFBB",X"FFD9",X"FFDC",X"FFCA",X"FFE5",X"0004",X"FFFA",X"FFDB",X"0012",X"0008",X"FFDA",X"FFDA",X"FFFE",X"000D",X"000E",X"002F",X"0020",X"FFE8",X"FFB6",X"FFAC",X"FFD7",X"FFF2",X"FFFB",X"0022",X"FFEA",X"FFB1",X"FFB6",X"FF9B",X"FF7B",X"FF99",X"FFE9",X"0002",X"0024",X"002A",X"FFF3",X"FFE4",X"FFF1",X"0011",X"000F",X"0015",X"FFFE",X"0007",X"0000",X"FFF6",X"FFEC",X"FFF6",X"FFF6",X"0005",X"FFF4",X"FFFC",X"003A",X"0078",X"0083",X"00A2",X"00C3",X"0098",X"0058",X"0050",X"0042",X"0029",X"004A",X"003E",X"0063",X"0065",X"0056",X"0061",X"0048",X"002B",X"0062",X"00B6",X"00E7",X"00D6",X"00D5",X"00BC",X"0088",X"0054",X"0042",X"001D",X"0010",X"0002",X"FFFE",X"FFFF",X"FFF3",X"FFB7",X"FF96",X"FF73",X"FF75",X"FF53",X"FF31",X"FF40",X"FF39",X"FF08",X"FF0C",X"FF2B",X"FF30",X"FF18",X"FF4B",X"FF8B",X"FF7C",X"FF69",X"FF58",X"FF1A",X"FF1B",X"FF3B",X"FF72",X"FF83",X"FFA5",X"FFAA",X"FF88",X"FF90",X"FFC7",X"FFB9",X"FFF5",X"006F",X"00A4",X"008C",X"0083",X"0065",X"0016",X"0007",X"0056",X"00A5",X"007E",X"005E",X"006E",X"0046",X"000E",X"0025",X"0032",X"0027",X"0010",X"002D",X"0039",X"000D",X"FFCC",X"FFC0",X"FFBB",X"FFAD",X"FFC6",X"FFD1",X"FFD5",X"FFCA",X"FFE4",X"FFEA",X"FFDF",X"FFA8",X"FFB3",X"FF9F",X"FFAE",X"FFB9",X"FFCB",X"FFD8",X"FFD6",X"FFB6",X"FF99",X"FF83",X"FF9D",X"FFD8",X"FFF2",X"0008",X"0005",X"FFD2",X"FF66",X"FF41",X"FF5B",X"FF89",X"FFA7",X"FFC6",X"FFCA",X"FFD8",X"FFC7",X"FFC0",X"FFA9",X"FF9A",X"FFAA",X"FFD0",X"FFFE",X"0006",X"FFE0",X"FFB9",X"FFB2",X"FFD7",X"0005",X"0018",X"FFEA",X"FFFA",X"001D",X"002B",X"0029",X"000B",X"0004",X"0024",X"0071",X"0089",X"0098",X"0087",X"0077",X"0069",X"0062",X"0087",X"009E",X"0092",X"009C",X"0099",X"0091",X"00BD",X"009B",X"0090",X"0068",X"007B",X"0081",X"007A",X"0066",X"0045",X"006A",X"007F",X"0076",X"004C",X"0034",X"0050",X"0057",X"0050",X"0004",X"FFF4",X"0040",X"006E",X"006D",X"0066",X"0069",X"005C",X"002B",X"FFF6",X"FFE3",X"FFD7",X"FFD7",X"FFF6",X"0027",X"0024",X"0014",X"0023",X"FFFF",X"002D",X"000E",X"FFF5",X"0022",X"FFFB",X"FFD5",X"FFCF",X"FFD3",X"FFA9",X"FF9C",X"FF9A",X"FF9F",X"FF8E",X"FF94",X"FF6F",X"FF57",X"FF3E",X"FF73",X"FF8F",X"FF80",X"FFC8",X"FFCD",X"FFD7",X"FFC9",X"FFCB",X"FF89",X"FF7A",X"FF9B",X"FFB5",X"FFBA",X"FF7F",X"FF8C",X"FF9B",X"FF7E",X"FF4D",X"FF56",X"FF59",X"FF7A",X"FFA9",X"FFF4",X"FFEB",X"FFA8",X"FFA7",X"FFAD",X"FFBD",X"FFDB",X"0019",X"0003",X"FFD1",X"FFBA",X"FFC4",X"FF92",X"FFB0",X"0015",X"002A",X"004A",X"006E",X"005B",X"0018",X"FFE6",X"FFE1",X"0019",X"004A",X"0074",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000");
begin
 
   
 process(resetN, CLK)
    variable num, curr_sound 		: integer;
	 type noteArrd is array (0 to 12) of integer;
	 variable dataTmp : noteArrd;
 begin

		if (resetN='0') then
			dataTmp := (others  => 0);
			num := 0;
			
		elsif(rising_edge(CLK)) then
			dataTmp := (others  => 0);
			num := 0;
			for i in 0 to 12 loop
				if conv_integer(addrArr(i)) > 0 then
					dataTmp(i) := conv_integer(sound0(conv_integer(addrArr(i))));--/num;
				end if;
			end loop;
		end if;
		Q <= conv_std_logic_vector(dataTmp(0) + dataTmp(1) + dataTmp(2) + dataTmp(3) + dataTmp(4) + dataTmp(5) + dataTmp(6) + dataTmp(7) + dataTmp(8) + dataTmp(9) + dataTmp(10) + dataTmp(11) + dataTmp(12), 16);
	end process;
	 

		   
end arch;