library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_signed.all ;
use ieee.std_logic_arith.all;
library work;
use work.pkg2.all;

entity sing_effect is
port(
  CLK     					: in std_logic;
  resetN 					: in std_logic;
  addrArr    				: in Arr_type;
  Q       					: out std_logic_vector(15 downto 0)
);
end sing_effect;

architecture arch of sing_effect is
	constant array_size 			: integer := 5000 ;
	
	signal Q_tmp       			:  std_logic_vector(15 downto 0) ;
	
	type table_type is array(0 to array_size - 1) of std_logic_vector(15 downto 0);
	constant sound0 : table_type := (X"003A",X"0014",X"FFCD",X"FFB9",X"FF84",X"FFA9",X"FFAD",X"FF7F",X"FF55",X"FF5F",X"FF60",X"FF60",X"FF4C",X"FF48",X"FF3E",X"FF6B",X"FF82",X"FF92",X"FF55",X"FF32",X"FF15",X"FF14",X"FF05",X"FF36",X"FF7E",X"FF9B",X"FF98",X"FF9F",X"FFA4",X"FF8F",X"FF9B",X"FF87",X"FFA4",X"FFCB",X"FFEC",X"000F",X"0010",X"FFF9",X"FFF5",X"0009",X"0032",X"003C",X"0032",X"002C",X"0048",X"0052",X"0069",X"009B",X"00AA",X"00A0",X"00CA",X"00F0",X"0128",X"014F",X"0125",X"00ED",X"00B3",X"00A6",X"00CC",X"00EA",X"00BC",X"009E",X"0087",X"006A",X"0065",X"0018",X"0007",X"0014",X"0021",X"0016",X"FFF9",X"FFBE",X"FF6E",X"FF40",X"FF4A",X"FF50",X"FF5A",X"FF68",X"FF91",X"FF8B",X"FF66",X"FF40",X"FF5D",X"FF9F",X"FFAF",X"FF9E",X"FF7E",X"FF80",X"FF8F",X"FFB0",X"FFA1",X"FF95",X"FFF3",X"0043",X"006B",X"004D",X"0030",X"005D",X"007A",X"008E",X"0097",X"009B",X"00AB",X"00BE",X"00CE",X"00D4",X"00C4",X"00BD",X"00AC",X"009E",X"009F",X"0052",X"0017",X"0012",X"0012",X"0008",X"FFEF",X"FFD9",X"FFEF",X"FFF9",X"FFFD",X"000D",X"000A",X"FFDE",X"FFB2",X"FF8B",X"FF89",X"FF99",X"FF77",X"FF4E",X"FF4F",X"FF63",X"FF5B",X"FF31",X"FF1D",X"FF4B",X"FF4E",X"FF4A",X"FF58",X"FF6C",X"FF8E",X"FFA4",X"FF8E",X"FF85",X"FF6C",X"FF64",X"FF81",X"FF8D",X"FF8F",X"FFAA",X"FFB9",X"FFB3",X"FF94",X"FF9C",X"FFB6",X"FFE4",X"FFFC",X"001A",X"001F",X"FFFE",X"0025",X"0025",X"001D",X"003F",X"0029",X"0026",X"005A",X"006D",X"004E",X"0022",X"FFF8",X"FFE3",X"FFEB",X"FFA6",X"FF75",X"FF7E",X"FFAA",X"FFB0",X"FF7A",X"FF63",X"FF74",X"FFB0",X"FFD0",X"FFC1",X"FFA9",X"FF98",X"FFAF",X"FFE8",X"FFE4",X"FFC0",X"FF9C",X"FF9B",X"FF9E",X"FFC3",X"FFD3",X"FFEB",X"0009",X"002A",X"001C",X"0007",X"0007",X"001C",X"0013",X"FFF5",X"001A",X"0043",X"0047",X"0069",X"0072",X"0062",X"008B",X"00AF",X"00CD",X"00D8",X"00E0",X"00FC",X"011E",X"00F9",X"00E1",X"00F7",X"00C7",X"009A",X"0092",X"0072",X"0064",X"005E",X"0027",X"0001",X"FFF0",X"FFCC",X"FF71",X"FF55",X"FF64",X"FF87",X"FFB5",X"FFC4",X"FFD4",X"FFDA",X"FFBC",X"FFB0",X"FF75",X"FF65",X"FF5E",X"FF6B",X"FFB2",X"FFBA",X"FF9A",X"FF7B",X"FF4F",X"FF4A",X"FF53",X"FF89",X"FFAA",X"FFD5",X"FFED",X"0003",X"0006",X"FFE6",X"0003",X"0019",X"0059",X"007E",X"008E",X"00A8",X"00B7",X"00A3",X"009C",X"00C1",X"00D8",X"00C6",X"00C0",X"00B3",X"0095",X"0079",X"008F",X"0072",X"005F",X"005D",X"004F",X"0075",X"007A",X"005C",X"0022",X"0016",X"0022",X"0030",X"FFE0",X"FF96",X"FFD1",X"FFD9",X"FFCA",X"FFB4",X"FFE5",X"001F",X"FFF6",X"FF97",X"FF48",X"FF56",X"FF7B",X"FF92",X"FF90",X"FF7C",X"FF6C",X"FF5F",X"FF68",X"FF6B",X"FF62",X"FF78",X"FF98",X"FF88",X"FF80",X"FF79",X"FF4F",X"FF4A",X"FF57",X"FF83",X"FFAC",X"FFF4",X"002D",X"004F",X"004E",X"0018",X"0012",X"0021",X"0014",X"000D",X"0011",X"004E",X"0052",X"0037",X"0039",X"0002",X"0004",X"000F",X"FFE7",X"FFFB",X"002B",X"003C",X"FFFD",X"FFB0",X"FF7E",X"FF9F",X"FFA9",X"FF89",X"FFA3",X"FFC7",X"FFE1",X"FFEE",X"FFE6",X"FFC7",X"FFC3",X"FFEE",X"FFE0",X"FFD0",X"FFBE",X"FFD6",X"FFBB",X"FF75",X"FF33",X"FF26",X"FF34",X"FF53",X"FF4D",X"FF47",X"FF49",X"FFA9",X"000F",X"0040",X"000D",X"0020",X"0025",X"001B",X"0049",X"004E",X"005C",X"0085",X"00AC",X"00DD",X"00BF",X"00AE",X"00A6",X"0081",X"0088",X"0096",X"00AD",X"00C7",X"0093",X"0086",X"0081",X"0050",X"0066",X"0076",X"0063",X"0093",X"008F",X"0073",X"006E",X"0050",X"0011",X"FFEE",X"FFE2",X"FFE3",X"FFE4",X"FFCE",X"FFCA",X"FFB6",X"FF90",X"FF7B",X"FF7C",X"FF49",X"FF3C",X"FF6C",X"FF80",X"FFA1",X"FFC2",X"FFCA",X"FFE7",X"FFF6",X"0002",X"0002",X"0012",X"0013",X"001B",X"FFF1",X"0005",X"0013",X"003D",X"005C",X"004A",X"005E",X"0047",X"0027",X"005A",X"0087",X"007D",X"0064",X"0059",X"002F",X"0005",X"0001",X"001D",X"0029",X"0042",X"009A",X"00C0",X"00A5",X"006A",X"0006",X"FFE3",X"FFF4",X"FFFF",X"0010",X"001D",X"0016",X"0017",X"FFF3",X"FF99",X"FF88",X"FFA3",X"FF7A",X"FF7B",X"FF55",X"FF30",X"FF11",X"FEE6",X"FEF7",X"FED9",X"FEB8",X"FEDE",X"FF1E",X"FF31",X"FF27",X"FEE1",X"FEA7",X"FE91",X"FE66",X"FE6D",X"FE88",X"FEB7",X"FEDD",X"FF12",X"FF58",X"FF5C",X"FF82",X"FF86",X"FFB3",X"FFF6",X"0007",X"0023",X"0011",X"002A",X"004A",X"0077",X"0084",X"00BE",X"0104",X"010C",X"011D",X"013F",X"0138",X"011E",X"00EE",X"00D3",X"00CD",X"00F2",X"00FD",X"0103",X"0118",X"00D5",X"00E1",X"00E1",X"00A9",X"0075",X"0047",X"0042",X"0034",X"0006",X"FFF8",X"FFFB",X"FFD9",X"FFCE",X"FFD3",X"FFDA",X"FFFF",X"001A",X"0017",X"003D",X"0011",X"FFE1",X"0010",X"FFF9",X"FFC0",X"FFCE",X"FFED",X"FFF8",X"FFE9",X"FFAB",X"FF73",X"FF56",X"FF5F",X"FF7E",X"FF7A",X"FF70",X"FF71",X"FF7D",X"FF71",X"FF8A",X"FFA6",X"FFDC",X"FFF5",X"000D",X"0002",X"FFF7",X"FFF8",X"0026",X"0025",X"001E",X"0059",X"00A8",X"00BD",X"00D1",X"0106",X"0148",X"015B",X"016F",X"019C",X"0194",X"0175",X"014B",X"011F",X"00F1",X"00DD",X"00A1",X"0055",X"0000",X"FFDF",X"FFC5",X"FF76",X"FF45",X"FF0D",X"FEFB",X"FED7",X"FE97",X"FE3A",X"FDFF",X"FDFE",X"FE04",X"FE0C",X"FDDE",X"FDDE",X"FDFE",X"FE45",X"FE87",X"FE6B",X"FEE3",X"FF67",X"0024",X"00B5",X"010C",X"018B",X"01CD",X"0204",X"01EB",X"01EE",X"0207",X"01EB",X"01CB",X"0185",X"00FC",X"0094",X"0054",X"FFF6",X"FF8D",X"FF5A",X"FF46",X"FF35",X"FEE5",X"FE62",X"FE42",X"FE09",X"FDC6",X"FD66",X"FCF8",X"FCB5",X"FCC5",X"FCBC",X"FCB8",X"FD28",X"FDEC",X"FECE",X"FFD2",X"00E9",X"024B",X"0395",X"04A2",X"051D",X"055B",X"05A9",X"0584",X"04F2",X"03FC",X"02F2",X"0208",X"0118",X"FFE9",X"FEC0",X"FDCD",X"FD10",X"FC7F",X"FC23",X"FBC7",X"FBA7",X"FB89",X"FB77",X"FB78",X"FB5C",X"FAF3",X"FB02",X"FAC4",X"FAF1",X"FBB8",X"FC9B",X"FE04",X"FF51",X"0153",X"035F",X"054E",X"075B",X"08DD",X"09D2",X"0A1B",X"0995",X"0877",X"0718",X"0612",X"0420",X"02C1",X"017E",X"FFF2",X"FF26",X"FE03",X"FD2A",X"FC4E",X"FC14",X"FC2E",X"FC29",X"FC5B",X"FC85",X"FCFD",X"FD07",X"FC98",X"FC0E",X"FB0D",X"FA6C",X"F98F",X"F97B",X"F9EF",X"FAA3",X"FC9B",X"FE50",X"011A",X"0386",X"05FE",X"0837",X"0972",X"0A3A",X"0A64",X"0931",X"0788",X"051C",X"03EC",X"0295",X"0149",X"002E",X"FEEC",X"FEB0",X"FE64",X"FDD2",X"FD60",X"FD05",X"FD0E",X"FD5F",X"FD39",X"FD1D",X"FD53",X"FD4E",X"FC93",X"FB40",X"FA02",X"F8D9",X"F808",X"F895",X"F913",X"F9F8",X"FBEA",X"FE76",X"0261",X"057B",X"094A",X"0AE3",X"0C84",X"0CFA",X"0C82",X"0ABD",X"072E",X"03CC",X"004B",X"FDF6",X"FDCB",X"FD0C",X"FC89",X"FDA6",X"FE89",X"FFBC",X"FF7C",X"FF1A",X"FF39",X"FF68",X"FF21",X"FDFD",X"FD1F",X"FC5C",X"FB6B",X"F9AF",X"F79F",X"F5D5",X"F4C4",X"F405",X"F52A",X"F5F9",X"F7C4",X"FA75",X"FE6A",X"0330",X"085B",X"0BD0",X"0E21",X"0FD0",X"1035",X"0FF4",X"0C69",X"0811",X"0343",X"003B",X"FEA8",X"FCDD",X"FCB0",X"FC60",X"FDF9",X"FF18",X"FF55",X"FFA8",X"FFB1",X"00BC",X"00C6",X"002C",X"FF37",X"FE5D",X"FD8E",X"FBD6",X"F965",X"F6CB",X"F505",X"F3AC",X"F366",X"F486",X"F5B6",X"F824",X"FB81",X"008E",X"0730",X"0C3A",X"0EEA",X"1135",X"11C5",X"1243",X"0F5E",X"0A82",X"04DE",X"00AA",X"FE9E",X"FC69",X"FA5D",X"F9AE",X"FA92",X"FCBF",X"FDD6",X"FE1D",X"FEBB",X"FFED",X"013A",X"012E",X"0014",X"FF52",X"FE98",X"FD06",X"FA86",X"F786",X"F530",X"F388",X"F24C",X"F308",X"F44E",X"F69B",X"F9DB",X"FF3B",X"066F",X"0C2A",X"100F",X"131D",X"1413",X"154C",X"12ED",X"0E90",X"08A9",X"03C8",X"0123",X"FE16",X"FB8E",X"F9D2",X"FA0A",X"FB9C",X"FC52",X"FC81",X"FCF9",X"FE7A",X"FFBB",X"FFB0",X"FF44",X"FE82",X"FD59",X"FBCD",X"F924",X"F620",X"F444",X"F19D",X"EFAB",X"EFD1",X"F1C5",X"F49B",X"F886",X"FD96",X"0495",X"0C54",X"10B0",X"14B6",X"155B",X"1625",X"149D",X"0FF1",X"09C8",X"0367",X"FF17",X"FC28",X"FB3B",X"F9CD",X"F9E1",X"FC02",X"FD29",X"FF76",X"FF2B",X"FF56",X"FFAC",X"002A",X"00AE",X"FF0E",X"FD92",X"FB82",X"F9A5",X"F7CA",X"F449",X"F107",X"EE9D",X"EE9C",X"F062",X"F1FC",X"F514",X"FAA6",X"0498",X"0C10",X"1200",X"154F",X"164F",X"186A",X"1699",X"12B0",X"0B33",X"04C4",X"00E4",X"FDB0",X"FAD6",X"F7F8",X"F6F9",X"F923",X"FB64",X"FC9B",X"FCAA",X"FDA0",X"FF17",X"0030",X"FFCB",X"FED6",X"FE92",X"FD1B",X"FAB1",X"F71F",X"F471",X"F0B3",X"EE00",X"EE80",X"F04A",X"F2F6",X"F6F6",X"FDEB",X"08B0",X"0EA1",X"1477",X"17F6",X"197E",X"1A6C",X"181E",X"1171",X"09CB",X"031F",X"FF3A",X"FBDB",X"F8DD",X"F746",X"F874",X"FB03",X"FCF9",X"FD8C",X"FE62",X"FF50",X"FFB4",X"004F",X"FF54",X"FDE3",X"FCD9",X"FA5B",X"F7A9",X"F378",X"F109",X"EDDB",X"EBEF",X"ED80",X"F051",X"F4BD",X"FBF5",X"0718",X"1034",X"166D",X"195F",X"1897",X"19C1",X"1678",X"10BD",X"0903",X"0130",X"FD7C",X"FAC4",X"F8A8",X"F7A3",X"F894",X"FC0B",X"FFD3",X"00F3",X"01A1",X"0359",X"02EE",X"022C",X"0069",X"FDC0",X"FCB5",X"FA29",X"F6EF",X"F371",X"EFEF",X"EE0B",X"ECF4",X"EE12",X"F397",X"F8AF",X"FE30",X"08B4",X"1392",X"16E1",X"19CB",X"15F4",X"1294",X"1111",X"08E3",X"FF7D",X"F883",X"F692",X"FAA3",X"FC66",X"FE81",X"0361",X"072A",X"09AD",X"0753",X"0107",X"FDA4",X"FBC1",X"F885",X"F7BF",X"F713",X"F8F3",X"F9E9",X"F778",X"F5B9",X"F007",X"EEB3",X"EAA0",X"EB52",X"F525",X"F8A0",X"0305",X"10EB",X"1C75",X"2156",X"1F40",X"1383",X"09FF",X"01E9",X"F76F",X"EF4B",X"EA84",X"F257",X"0309",X"0B5B",X"1446",X"169E",X"145E",X"10B1",X"0245",X"F494",X"EF3F",X"ECEF",X"F1B1",X"F7B8",X"FB20",X"00DE",X"0231",X"FDF6",X"F977",X"EE32",X"E9E1",X"E4E8",X"E02D",X"EE2E",X"F7D0",X"04C9",X"19CE",X"2799",X"27D3",X"2217",X"0E31",X"FECD",X"F5DA",X"EB6E",X"E820",X"EC8D",X"FCA4",X"1216",X"1AEB",X"1E35",X"187A",X"0D07",X"024C",X"F23C",X"E96D",X"ECED",X"F489",X"FF2B",X"058B",X"06D2",X"0706",X"01DD",X"F841",X"F1D2",X"E9DC",X"E839",X"E5EA",X"E7CA",X"F7EB",X"0599",X"13CA",X"27AB",X"2609",X"1CD8",X"10E6",X"FB89",X"EF9E",X"EB78",X"E588",X"F02D",X"FED6",X"13EA",X"2245",X"2227",X"18D4",X"0ACC",X"F9FE",X"ED9F",X"E559",X"E97B",X"F79B",X"0374",X"09F5",X"09FF",X"0639",X"0045",X"F7D1",X"EF15",X"EB21",X"E83C",X"E6A4",X"E5F5",X"F2BD",X"03F2",X"1377",X"228C",X"2799",X"1C01",X"10A2",X"FE2B",X"ED8D",X"E996",X"E861",X"F0E2",X"0019",X"159A",X"23B1",X"2369",X"179A",X"074E",X"F6DD",X"ECCA",X"E696",X"EC13",X"FA38",X"06FF",X"0B94",X"095F",X"0360",X"FD4E",X"F5FC",X"EE4B",X"EB05",X"EB23",X"EB55",X"E69C",X"F03A",X"0414",X"1162",X"1D9A",X"26E2",X"1B84",X"0FD8",X"FE50",X"ED07",X"E907",X"EA76",X"F0C0",X"006D",X"14AE",X"23BD",X"2342",X"1650",X"0516",X"F422",X"EBD6",X"E823",X"EE45",X"FCA0",X"0924",X"0D2C",X"0874",X"018D",X"FC15",X"F49E",X"EF52",X"EC7B",X"EB6A",X"ED6C",X"E9FD",X"EF1D",X"023B",X"0D53",X"1958",X"285D",X"1E0A",X"0FDA",X"00E2",X"EF18",X"E9A9",X"EC2F",X"EFC5",X"FF47",X"1514",X"2326",X"22B4",X"1542",X"038C",X"F416",X"EC34",X"E949",X"EFDA",X"FCE4",X"0903",X"0C72",X"071D",X"FFCE",X"FA35",X"F530",X"F002",X"EEB7",X"ED76",X"EB1A",X"E6AB",X"ECCA",X"028B",X"11D7",X"1E33",X"2B26",X"2004",X"10C1",X"FFE6",X"ECA8",X"E755",X"EB09",X"F234",X"0437",X"1999",X"265C",X"248F",X"1470",X"007C",X"EFBA",X"E8ED",X"E8C2",X"F2DB",X"00CD",X"0C79",X"0EBE",X"0710",X"FEC2",X"F8B1",X"F3C8",X"EFA8",X"ED6E",X"EBEE",X"EBDB",X"E70B",X"EF88",X"046C",X"13FB",X"2347",X"2AE4",X"1B90",X"0CF8",X"FA67",X"E92B",X"E6DB",X"EA35",X"F4E7",X"08D7",X"1D3C",X"27A3",X"2204",X"0E2E",X"FA2B",X"EAAF",X"E64E",X"EA85",X"F67D",X"0455",X"0EE3",X"0EFD",X"050D",X"FBE6",X"F502",X"F131",X"EDC4",X"EE4C",X"ECE3",X"E99E",X"E434",X"F2B6",X"094C",X"1A04",X"2A0E",X"2928",X"15B2",X"080A",X"F4C4",X"E627",X"E773",X"EC32",X"FB0D",X"10B7",X"232A",X"28C1",X"1EB0",X"089C",X"F361",X"E71D",X"E5DD",X"EDFB",X"FB57",X"08E6",X"0F8D",X"0C73",X"003D",X"F92C",X"F436",X"F165",X"EDFC",X"EBF0",X"EA12",X"E6FE",X"E59A",X"F8FC",X"0E4C",X"1F30",X"2E07",X"249C",X"0F9F",X"FF82",X"ED03",X"E38B",X"E791",X"EFA6",X"023A",X"197D",X"289C",X"2789",X"1859",X"FFC3",X"ECC2",X"E6E1",X"E7F9",X"F39B",X"01CF",X"0BED",X"0F47",X"08AA",X"FCE4",X"F861",X"F50F",X"F314",X"F1BF",X"EE0C",X"EA4F",X"E419",X"E833",X"FE54",X"12CE",X"22E5",X"2E43",X"1F10",X"0CBA",X"F9EA",X"E80E",X"E50B",X"EA75",X"F418",X"089D",X"1EDE",X"29E4",X"251E",X"10A7",X"F84C",X"E94C",X"E5C0",X"EB35",X"F90C",X"055F",X"0DB4",X"0D6A",X"02E2",X"FA8A",X"F715",X"F4B0",X"F336",X"F09A",X"EC80",X"E8A9",X"E1E4",X"EF52",X"0641",X"18DF",X"29F7",X"2AE0",X"15FE",X"05D1",X"F1C7",X"E419",X"E70E",X"EE3F",X"FC0E",X"1312",X"2585",X"298F",X"1FB0",X"0776",X"F15F",X"E886",X"E8B9",X"F319",X"018F",X"0A4B",X"0EF4",X"0B47",X"FEB6",X"F94B",X"F655",X"F44F",X"F316",X"EFA1",X"ED23",X"E914",X"E4B3",X"F5D2",X"0B07",X"1BDB",X"2D28",X"25F5",X"0EE6",X"FDC9",X"EBE4",X"E388",X"E88D",X"EFB7",X"FFE1",X"1780",X"26E4",X"26C4",X"1848",X"FEC5",X"EBFF",X"E6B2",X"EA83",X"F777",X"0382",X"0AFB",X"0CD3",X"0505",X"FA83",X"F60C",X"F3DD",X"F3BF",X"F313",X"F02F",X"ECD3",X"E625",X"E838",X"FB39",X"0FE6",X"21B6",X"2DC7",X"20A7",X"0C99",X"F905",X"E88F",X"E499",X"EA32",X"F46F",X"08F0",X"1F20",X"295A",X"246D",X"0FAB",X"F722",X"E980",X"E869",X"F09D",X"FEAC",X"088C",X"0D6F",X"0B5D",X"0138",X"F8F6",X"F5A0",X"F4CB",X"F4EB",X"F39F",X"EEDE",X"EA12",X"E394",X"EDE8",X"032D",X"1720",X"2660",X"294B",X"177D",X"061E",X"F1BD",X"E400",X"E500",X"EC45",X"F903",X"1020",X"227C",X"270C",X"1DE9",X"0645",X"F0C0",X"E85C",X"E999",X"F4BC",X"019E",X"08F1",X"0BA6",X"0692",X"FCA6",X"F894",X"F691",X"F71C",X"F614",X"F30B",X"EDE8",X"E80D",X"E4A4",X"F4A2",X"09DF",X"1E08",X"2D85",X"2944",X"1400",X"00C1",X"ED4C",X"E3FD",X"E776",X"EFE7",X"FFDE",X"16FF",X"26F2",X"2799",X"17EB",X"0010",X"ED7F",X"E7E1",X"ED74",X"FA6E",X"046D",X"0A86",X"09E7",X"024D",X"FAAB",X"F854",X"F72B",X"F767",X"F476",X"EFBF",X"E9B6",X"E4B2",X"E8EE",X"FB72",X"0F92",X"2227",X"2C9B",X"2090",X"0CE7",X"F74F",X"E68D",X"E40D",X"E9E0",X"F4BD",X"08F5",X"1CC3",X"2563",X"2121",X"0DB1",X"F76A",X"EB6C",X"EA5E",X"F290",X"FEC4",X"0634",X"0975",X"0759",X"0054",X"FBA7",X"FA07",X"F885",X"F694",X"F348",X"ED45",X"E815",X"E405",X"F184",X"05CF",X"1995",X"2A4C",X"2A77",X"1758",X"0561",X"F022",X"E47C",X"E6B3",X"EE06",X"FBB0",X"1194",X"2210",X"258F",X"1B05",X"046D",X"F081",X"E8F8",X"EBFD",X"F6D3",X"014E",X"076D",X"0830",X"03B5",X"FC81",X"F9F2",X"F838",X"F69F",X"F465",X"F0C2",X"E9C3",X"E4FF",X"E649",X"F68B",X"0A49",X"1D83",X"2C16",X"24B0",X"10BE",X"FCE5",X"EB05",X"E564",X"EA1A",X"F308",X"03BC",X"1734",X"23D2",X"22FF",X"12C1",X"FCF5",X"ED98",X"E999",X"F0E1",X"FCF0",X"0537",X"0990",X"07D2",X"0143",X"FBAB",X"F9D5",X"F97F",X"F770",X"F4A9",X"F052",X"EA1E",X"E56A",X"EF26",X"FFB0",X"1109",X"2158",X"2977",X"1D3B",X"0B5B",X"F5EF",X"E7E8",X"E769",X"EE23",X"F83F",X"0A1C",X"1A45",X"222C",X"1D1D",X"0AB0",X"F63A",X"EBC8",X"EC4F",X"F537",X"FFEA",X"066F",X"07F2",X"04E6",X"FDD3",X"FA94",X"F9A7",X"F867",X"F590",X"F2F2",X"EC8D",X"E85D",X"E63D",X"F269",X"049D",X"17D2",X"25FC",X"2725",X"166D",X"0572",X"F1FA",X"E77A",X"E982",X"F1BE",X"FDF6",X"117D",X"1FE1",X"2329",X"1904",X"04AA",X"F20B",X"EBCD",X"EFDA",X"FAAB",X"0434",X"090C",X"08CF",X"03FD",X"FCFB",X"FAB0",X"F9B9",X"F91E",X"F710",X"F387",X"ECAF",X"E8EF",X"E8EA",X"F5FF",X"06DD",X"1940",X"278B",X"23F8",X"1212",X"0061",X"EDF6",X"E6E6",X"EAFE",X"F355",X"01F3",X"144A",X"1F34",X"1FBA",X"11E7",X"FC97",X"ED9E",X"E969",X"EFDB",X"FC2E",X"0403",X"07C3",X"05CF",X"FF71",X"FAB3",X"F949",X"F86E",X"F762",X"F4FA",X"F041",X"E981",X"E591",X"EC97",X"FCCC",X"0CD7",X"1D15",X"278B",X"209E",X"0EED",X"FC0D",X"EC39",X"E85B",X"EE6F",X"F891",X"09C2",X"1ACE",X"217A",X"1DA9",X"0D36",X"F8FF",X"EE91",X"EDC9",X"F554",X"FF9A",X"055C",X"06E8",X"03D3",X"FDB7",X"FAF9",X"F950",X"F7AA",X"F639",X"F3CA",X"EF74",X"EB28",X"E68B",X"EE7F",X"FEF7",X"0EF7",X"1D6D",X"25C2",X"1B6A",X"0A20",X"F78E",X"EA7D",X"E8EF",X"EF20",X"F85E",X"0A2A",X"1962",X"1F19",X"1A48",X"08B6",X"F6C1",X"EE5B",X"EE3A",X"F6C0",X"FFF1",X"04EF",X"06E5",X"0339",X"FD0F",X"FAC3",X"F9A8",X"F948",X"F6F2",X"F439",X"EFAD",X"EC10",X"E9EB",X"F381",X"02AB",X"1362",X"1F61",X"2562",X"1AA0",X"0900",X"F5C0",X"EA8B",X"EA68",X"F24F",X"FCBB",X"0EE3",X"1C0D",X"2138",X"1916",X"05B6",X"F4FE",X"EEB8",X"F09F",X"F9D4",X"01C8",X"064E",X"0671",X"026E",X"FCFA",X"FA78",X"F857",X"F7F6",X"F5A4",X"F336",X"EEA5",X"EB00",X"E912",X"F3FB",X"03F4",X"143D",X"1F5D",X"21BD",X"153F",X"0602",X"F3C2",X"EA58",X"EB83",X"F2FD",X"FEB3",X"1105",X"1C54",X"1E57",X"1461",X"0267",X"F415",X"EF15",X"F1AA",X"FB4B",X"026C",X"0618",X"060B",X"017A",X"FC9E",X"FAE9",X"F941",X"F921",X"F6BB",X"F400",X"F036",X"EBE4",X"EA51",X"F563",X"04AB",X"14EE",X"1FAC",X"2104",X"15CC",X"0588",X"F3E1",X"EB57",X"EC5C",X"F388",X"FF7E",X"10B0",X"1C67",X"1E7C",X"1447",X"01A1",X"F2AD",X"ED92",X"F07E",X"F9CC",X"0180",X"0591",X"05DF",X"0147",X"FBFC",X"FA05",X"F83A",X"F78C",X"F499",X"F151",X"ECD8",X"E833",X"E7E5",X"F421",X"0485",X"1517",X"2036",X"2195",X"1677",X"05BC",X"F305",X"E96D",X"EAEB",X"F339",X"00A3",X"12F3",X"1DC0",X"1E9C",X"13DA",X"004D",X"F28C",X"EE6B",X"F19F",X"FB1A",X"01B1",X"0568",X"0590",X"0116",X"FD40",X"FB88",X"F9B3",X"F8C6",X"F5D4",X"F26D",X"EE04",X"E8AB",X"E938",X"F62C",X"0711",X"161D",X"1FBA",X"2104",X"1656",X"05A9",X"F3C3",X"EA51",X"EBF9",X"F423",X"01B1",X"139E",X"1DE7",X"1E68",X"12CE",X"0032",X"F3ED",X"EFAF",X"F2E0",X"FC20",X"021A",X"05C7",X"0655",X"01A0",X"FD9F",X"FBA4",X"F9F7",X"F934",X"F601",X"F221",X"ED65",X"E883",X"E969",X"F67C",X"07B4",X"1633",X"1F18",X"202C",X"158D",X"05A5",X"F4DE",X"EB0D",X"EC64",X"F4FC",X"02A9",X"14BF",X"1EE6",X"1E98",X"130F",X"0054",X"F3C1",X"F00D",X"F2C0",X"FBD9",X"021F",X"05B4",X"0687",X"0255",X"FDD4",X"FB77",X"F8D3",X"F77D",X"F413",X"F0DE",X"EDEB",X"EA76",X"EB5A",X"F6C8",X"064D",X"1421",X"1B8D",X"1CD5",X"144D",X"0479",X"F49D",X"EC44",X"ED12",X"F58A",X"0323",X"13E3",X"1CAE",X"1C55",X"0FD4",X"FDBD",X"F352",X"F03C",X"F363",X"FCD4",X"02DD",X"0603",X"0615",X"0139",X"FCAF",X"F9C9",X"F812",X"F750",X"F401",X"F17E",X"EE4C",X"EA54",X"EB66",X"F71B",X"05B9",X"12C1",X"1B26",X"1BCD",X"12C7",X"04D6",X"F585",X"ED73",X"EF25",X"F6C7",X"03A6",X"132C",X"1B5F",X"1B3D",X"0E95",X"FD6C",X"F36B",X"F03A",X"F490",X"FDF3",X"038A",X"06F1",X"0633",X"0007",X"FA3C",X"F738",X"F65D",X"F6C9",X"F497",X"F17D",X"ECB6",X"E90E",X"EC9C",X"F96A",X"07C3",X"14BE",X"1C5D",X"1C30",X"137B",X"04CD",X"F452",X"EC08",X"EE05",X"F70C",X"05DD",X"163C",X"1C6A",X"1ABE",X"0D4D",X"FB6F",X"F210",X"F02E",X"F590",X"FEC3",X"03E7",X"0743",X"05AF",X"FFA1",X"FB14",X"F819",X"F74F",X"F795",X"F47A",X"F1FD",X"EDF8",X"E9E3",X"EDB5",X"F90E",X"071A",X"154F",X"1CAE",X"1D18",X"1511",X"05A0",X"F675",X"EE77",X"EF65",X"F832",X"068B",X"165B",X"1DC9",X"1B5F",X"0DCC",X"FCC5",X"F2FE",X"F1B2",X"F6BE",X"FF04",X"03E6",X"0634",X"049B",X"FF3B",X"FA9D",X"F7BD",X"F76F",X"F7C1",X"F5C9",X"F29F",X"ED9D",X"E955",X"EE51",X"FA04",X"07BE",X"1437",X"1C37",X"1C94",X"1496",X"04E5",X"F51C",X"EC77",X"EE44",X"F708",X"06B2",X"1640",X"1C98",X"1AD6",X"0D19",X"FB62",X"F247",X"F056",X"F5EA",X"FE43",X"02CB",X"05ED",X"0452",X"FECD",X"FA9A",X"F779",X"F731",X"F662",X"F486",X"F2D7",X"EDD2",X"E948",X"EDA4",X"F95D",X"06DF",X"1350",X"1CC1",X"1CF1",X"13B8",X"04A9",X"F4A7",X"EC60",X"EF06",X"F721",X"06F8",X"1689",X"1BD9",X"198C",X"0BDB",X"FAEE",X"F2C1",X"F16E",X"F740",X"FEE3",X"02DD",X"04FE",X"02A5",X"FD87",X"FA0C",X"F762",X"F753",X"F6F6",X"F420",X"F19D",X"ED3E",X"E9D0",X"F002",X"FC2E",X"08D4",X"1528",X"1CF7",X"1BDF",X"1294",X"02C0",X"F3D7",X"ED3C",X"F047",X"F968",X"093B",X"183D",X"1D1B",X"1843",X"0A01",X"F93E",X"F07B",X"F0EA",X"F7C2",X"FF8D",X"0436",X"05AC",X"0344",X"FDDA",X"F960",X"F757",X"F765",X"F633",X"F407",X"F0BA",X"ED00",X"EB39",X"F0F6",X"FCCF",X"08FF",X"1480",X"1CD8",X"1B7F",X"122A",X"0308",X"F44F",X"EE53",X"F1D0",X"FAE1",X"0B6F",X"187E",X"1BD7",X"1702",X"08E7",X"FA5C",X"F305",X"F2E6",X"F9B3",X"FFA6",X"0318",X"04A8",X"0222",X"FE00",X"FAD8",X"F8F2",X"F8C2",X"F67B",X"F3B5",X"F0C1",X"ECC3",X"EB72",X"F157",X"FD9C",X"0A3C",X"1520",X"1C5A",X"1A7D",X"10FE",X"0228",X"F47F",X"EF0F",X"F236",X"FB12",X"0B54",X"1962",X"1CEF",X"1658",X"0785",X"F8EA",X"F196",X"F1F5",X"F8AA",X"FF03",X"02D7",X"03C1",X"011A",X"FCD9",X"F98F",X"F81F",X"F845",X"F6DB",X"F482",X"F091",X"ED07",X"EB2F",X"F07C",X"FD59",X"0A9E",X"15D2",X"1DBD",X"1AF4",X"104E",X"00F2",X"F2F0",X"EE3E",X"F26D",X"FC64",X"0D89",X"197E",X"1BB5",X"14B1",X"055D",X"F86E",X"F2C4",X"F374",X"FA97",X"0000",X"0315",X"0391",X"0016",X"FBFF",X"F9A3",X"F8A8",X"F871",X"F5D8",X"F309",X"EF11",X"EBBF",X"EA70",X"F0EC",X"FE45",X"0B99",X"1653",X"1CCE",X"195E",X"0E21",X"FEC0",X"F1D9",X"EDD7",X"F2C7",X"FD60",X"0E11",X"1946",X"1B3F",X"1315",X"038D",X"F7C4",X"F2F5",X"F3D9",X"FAC3",X"FF90",X"0271",X"02D5",X"FF47",X"FB8F",X"F96E",X"F87D",X"F83B",X"F639",X"F359",X"EF53",X"EBB5",X"EA9A",X"F3AF",X"01F4",X"0DF9",X"185F",X"1D18",X"176F",X"0BD4",X"FCEF",X"F1CC",X"EFC0",X"F51D",X"0110",X"1097",X"1993",X"1A21",X"1089",X"015B",X"F70C",X"F3CE",X"F69E",X"FCD4",X"00D9",X"02BA",X"01B0",X"FF00",X"FC08",X"FA86",X"FA36",X"F87F",X"F590",X"F233",X"ED99",X"EB7F",X"EC9A",X"F65C",X"055D",X"1190",X"19F1",X"1BF4",X"146A",X"0776",X"F9A1",X"F114",X"F144",X"F786",X"05A5",X"141E",X"199F",X"188B",X"0D74",X"FE6B",X"F68B",X"F46E",X"F8BC",X"FE6B",X"00FA",X"02C9",X"0163",X"FDBA",X"FAE8",X"F975",X"F9D0",X"F8E7",X"F545",X"F11F",X"EDD8",X"EBC2",X"EEFE",X"FADC",X"07C6",X"129E",X"1AE1",X"1A6D",X"11C7",X"03BC",X"F5D4",X"EF5D",X"F14B",X"F936",X"093E",X"16AE",X"1A76",X"14B7",X"07D0",X"FAFA",X"F4CB",X"F573",X"FB19",X"FFC1",X"0233",X"0298",X"004A",X"FD18",X"FA99",X"F9AA",X"F8CF",X"F784",X"F544",X"F0AD",X"ED01",X"EB80",X"F204",X"FF11",X"0BEB",X"15EC",X"1BAB",X"1759",X"0C91",X"FE13",X"F247",X"EEE3",X"F347",X"FEE9",X"0EEF",X"1836",X"19A3",X"101F",X"010E",X"F79E",X"F39E",X"F622",X"FCC6",X"0092",X"02DC",X"0231",X"FECD",X"FBED",X"FA5C",X"FA00",X"F8BD",X"F645",X"F3C8",X"EFE0",X"EC87",X"ED72",X"F6E9",X"0467",X"1025",X"189F",X"1A76",X"13B1",X"06F9",X"F924",X"F03E",X"EF99",X"F604",X"052B",X"1373",X"18F8",X"1640",X"0A67",X"FB9A",X"F467",X"F3FB",X"F8CD",X"FE81",X"0172",X"023E",X"00C0",X"FDB7",X"FAD9",X"FA1D",X"F9C4",X"F741",X"F4B3",X"F160",X"EE75",X"EBDA",X"F013",X"FC47",X"0994",X"1451",X"1B8E",X"193A",X"0FE9",X"0186",X"F536",X"F022",X"F359",X"FCD6",X"0C9A",X"17C6",X"19BA",X"1219",X"0437",X"F990",X"F5C5",X"F710",X"FC8F",X"0037",X"0156",X"005F",X"FDEC",X"FB28",X"FA75",X"FB21",X"FB1D",X"F7BD",X"F39E",X"EF16",X"EB7A",X"EBDD",X"F48F",X"023C",X"0F66",X"18B7",X"1C34",X"16D0",X"0ACA",X"FC6B",X"F260",X"F071",X"F5D4",X"033E",X"1218",X"18D2",X"17CD",X"0D58",X"FEF6",X"F714",X"F56C",X"F90B",X"FE33",X"00D3",X"0168",X"FFDC",X"FCDD",X"FB03",X"FB32",X"FC17",X"FA22",X"F60C",X"F18A",X"ED59",X"EB15",X"EEBA",X"FA33",X"074A",X"126D",X"1AFB",X"1AC7",X"126F",X"046F",X"F641",X"EFCF",X"F27B",X"FAE5",X"0AD9",X"16FA",X"1975",X"1296",X"0568",X"FA70",X"F5C5",X"F673",X"FBE5",X"FF54",X"008D",X"0022",X"FD1F",X"FA76",X"F9FF",X"FA94",X"FA54",X"F77D",X"F3DE",X"EF28",X"EB14",X"EABF",X"F2FA",X"00BD",X"0E2A",X"17EE",X"1BDC",X"16C2",X"0AFD",X"FC5D",X"F201",X"F00C",X"F566",X"028D",X"1168",X"182A",X"179E",X"0DAD",X"FEF4",X"F71A",X"F629",X"F97F",X"FE4B",X"FFE9",X"FFD8",X"FE5A",X"FBD4",X"FAAA",X"FAF7",X"FB86",X"F96D",X"F51F",X"F0C7",X"EBBE",X"E928",X"EE16",X"F9C4",X"0746",X"128A",X"1AEB",X"1AD4",X"120D",X"0402",X"F67C",X"EFF5",X"F20D",X"FA97",X"0AA7",X"16E2",X"1960",X"12AF",X"05EF",X"FB6D",X"F707",X"F7B7",X"FD02",X"0040",X"00C3",X"0058",X"FDAF",X"FBAE",X"FBB3",X"FC6B",X"FC5B",X"F8B0",X"F429",X"EE8B",X"EB45",X"EB8B",X"F335",X"00A4",X"0D57",X"16C7",X"1BD9",X"174C",X"0BDC",X"FD29",X"F280",X"F075",X"F5FD",X"039E",X"1257",X"1769",X"1590",X"0C10",X"FF45",X"F8B5",X"F7D6",X"FACD",X"FEAC",X"FFF8",X"FFB5",X"FDF9",X"FBEF",X"FB0F",X"FB9D",X"FD1F",X"FB59",X"F694",X"F283",X"EDD4",X"EB02",X"EF0F",X"F9B5",X"0696",X"1216",X"19F1",X"19B1",X"11BB",X"03B7",X"F70E",X"F137",X"F31A",X"FB5A",X"0A58",X"1567",X"17F1",X"108B",X"044E",X"FB98",X"F7F7",X"F98D",X"FEC4",X"0111",X"00D8",X"FF18",X"FBE0",X"FA67",X"FB17",X"FCD2",X"FD1F",X"F951",X"F502",X"EFEF",X"EC38",X"EBF7",X"F39D",X"001D",X"0CD4",X"158D",X"19EA",X"15C2",X"0AD5",X"FCC4",X"F346",X"F197",X"F71A",X"0435",X"1124",X"1516",X"128A",X"096A",X"FE24",X"F87E",X"F7E4",X"FB94",X"FF48",X"FF9F",X"FECB",X"FCD3",X"FB01",X"FA5C",X"FB4A",X"FC96",X"FB02",X"F6AC",X"F259",X"ED81",X"EB66",X"F03E",X"FAB1",X"05D9",X"0FFE",X"16D9",X"1755",X"104E",X"0371",X"F7B3",X"F287",X"F40E",X"FC5D",X"0B10",X"13F4",X"154A",X"0D56",X"0174",X"FA9F",X"F805",X"F98F",X"FE9A",X"0014",X"0038",X"FECC",X"FBC4",X"FAB0",X"FB0E",X"FC87",X"FCBC",X"F91F",X"F4F0",X"F126",X"ED91",X"ECD3",X"F462",X"00ED",X"0D08",X"1525",X"18EF",X"14B3",X"0A89",X"FD76",X"F4D5",X"F344",X"F84C",X"054F",X"1187",X"1436",X"10E6",X"06E0",X"FCB1",X"F8AD",X"F8BF",X"FCEE",X"00AD",X"00CF",X"FF8F",X"FCE6",X"FA9F",X"FA80",X"FC27",X"FDC7",X"FB94",X"F727",X"F398",X"EEF1",X"ECD3",X"F231",X"FC0B",X"06C0",X"1190",X"1861",X"17A0",X"1014",X"03F0",X"F964",X"F465",X"F5F3",X"FE07",X"0C2F",X"14BE",X"1513",X"0D45",X"01D0",X"FB04",X"F970",X"FB10",X"0009",X"015B",X"008C",X"FEFE",X"FBCB",X"FA5A",X"FB18",X"FC6D",X"FC5F",X"F92F",X"F4ED",X"F029",X"ECE2",X"EC5A",X"F3EC",X"00AD",X"0BF7",X"1423",X"1878",X"1486",X"0B60",X"FEE8",X"F5EE",X"F3AF",X"F7A2",X"02D6",X"0FD1",X"13DD",X"1255",X"08DF",X"FD6F",X"F976",X"F965",X"FBEE",X"FF42",X"FF10",X"FE5F",X"FC74",X"FA37",X"FA54",X"FBB5",X"FCBA",X"FB00",X"F615",X"F22B",X"EEA8",X"EC0C",X"EE6C",X"F7C9",X"03A2",X"0E9D",X"164A",X"1763",X"1149",X"06AE",X"FB92",X"F520",X"F565",X"FA7F",X"0788",X"1293",X"1439",X"0F20",X"0521",X"FC1C",X"F991",X"FA31",X"FE10",X"FFF5",X"FEE0",X"FE0D",X"FC5A",X"FB19",X"FBFD",X"FD1C",X"FD41",X"FA04",X"F50A",X"F108",X"EEAF",X"ED87",X"F118",X"FAE3",X"063E",X"109C",X"180C",X"16EC",X"0FA3",X"03E9",X"F9DA",X"F59D",X"F741",X"FE2F",X"0B4E",X"1345",X"1430",X"0CE9",X"023F",X"FC45",X"FAD2",X"FBDB",X"FF36",X"FF86",X"FE6F",X"FCD2",X"FA99",X"FAA9",X"FBBA",X"FCE4",X"FBA7",X"F7D3",X"F3CB",X"F071",X"EEE0",X"EE0F",X"F2C8",X"FE63",X"0955",X"11C3",X"1730",X"1452",X"0CC8",X"01BE",X"F95A",X"F6BB",X"F8E0",X"0107",X"0CDC",X"1157",X"1237",X"0AB3",X"FFED",X"FCC5",X"FC97",X"FE34",X"0118",X"0030",X"FEC1",X"FD2B",X"FAD7",X"FB58",X"FCB2",X"FDC2",X"FC4E",X"F7DA",X"F3CF",X"F089",X"EE68",X"EEAC",X"F519",X"0136",X"0BA3",X"131E",X"16DA",X"134E",X"0B57",X"00B9",X"F99B",X"F839",X"FAAC",X"03C8",X"0E83",X"121A",X"10AE",X"0812",X"FDC8",X"FB39",X"FB0A",X"FD22",X"FFC6",X"FEF9",X"FDC3",X"FC70",X"FA65",X"FAFF",X"FC19",X"FC91",X"FA7F",X"F680",X"F319",X"F0C0",X"EDD4",X"ED45",X"F5B2",X"018C",X"0BB0",X"1465",X"15D0",X"10CE",X"08B4",X"FE52",X"F80F",X"F78E",X"FA36",X"04E3",X"0F7D",X"125E",X"0F3D",X"0663",X"FD4E",X"FAD8",X"FB30",X"FE16",X"FF38",X"FDFA",X"FCE7",X"FB7E",X"FA75",X"FB18",X"FC51",X"FC79",X"F9A6",X"F5BB",X"F2B6",X"EFAD",X"EE09",X"EF5D",X"F7D6",X"0374",X"0D54",X"14B1",X"14C9",X"0EF8",X"0656",X"FD85",X"F849",X"F8FF",X"FD1C",X"0868",X"10D5",X"1200",X"0D6F",X"0477",X"FDC1",X"FC7A",X"FCBD",X"FF73",X"FFB0",X"FDE2",X"FC8F",X"FAFC",X"FAF0",X"FC1A",X"FD32",X"FC87",X"F914",X"F5A5",X"F2A4",X"EFF1",X"EE8D",X"F0BD",X"FA25",X"0572",X"0F85",X"168D",X"147F",X"0DD1",X"046F",X"FBC9",X"F888",X"F98C",X"FDE7",X"0949",X"10CF",X"11F5",X"0C5C",X"02A1",X"FCB4",X"FBC1",X"FC96",X"FFDF",X"FFB6",X"FE2C",X"FCD7",X"FB3B",X"FB96",X"FCEB",X"FD77",X"FC80",X"F8E3",X"F4B1",X"F123",X"EFF5",X"EF4C",X"F333",X"FD6C",X"07D6",X"0FD5",X"14E5",X"1289",X"0C3A",X"0332",X"FC38",X"F9EA",X"FB2E",X"009A",X"0B9D",X"11BD",X"11E6",X"0B5B",X"0223",X"FDB0",X"FCF8",X"FDCC",X"FFF3",X"FF43",X"FE28",X"FD4A",X"FC49",X"FC94",X"FD74",X"FD55",X"FB26",X"F70F",X"F3B5",X"F10A",X"F005",X"EF80",X"F4EB",X"FE65",X"08BF",X"10B7",X"1424",X"10D1",X"0A5F",X"00B0",X"FB12",X"F9DC",X"FB33",X"01AD",X"0BF2",X"10A3",X"104D",X"08F2",X"FFF6",X"FCB5",X"FCBA",X"FE98",X"0047",X"FE88",X"FD49",X"FC02",X"FB4D",X"FC6D",X"FD34",X"FCBE",X"FA43",X"F5A0",X"F2BF",X"F0CC",X"EF79",X"EF17",X"F594",X"FFCC",X"0993",X"0FD0",X"11E0",X"0E36",X"0810",X"FFBA",X"FAF7",X"F9E4",X"FB87",X"0266",X"0BF0",X"0FFE",X"0EB2",X"07B6",X"FF7D",X"FC86",X"FCBE",X"FEC4",X"FFD5",X"FE81",X"FD46",X"FC70",X"FC20",X"FD19",X"FE19",X"FD47",X"FA11",X"F589",X"F254",X"F085",X"EFCD",X"F051",X"F770",X"0160",X"0ACB",X"1179",X"12A3",X"0EDE",X"081E",X"FF49",X"FB13",X"FA85",X"FC6D",X"04D0",X"0D59",X"0FE4",X"0DC6",X"05FA",X"FF43",X"FDE7",X"FD68",X"FF3E",X"FFC7",X"FDF5",X"FD6B",X"FCC4",X"FCD0",X"FE2B",X"FE97",X"FD76",X"FA24",X"F5B2",X"F319",X"F165",X"F0B0",X"F206",X"F8D5",X"0276",X"0B33",X"1043",X"10B2",X"0D45",X"0745",X"FFD8",X"FC11",X"FB93",X"FD76",X"0595",X"0D9E",X"0FFD",X"0CB5",X"0566",X"FF80",X"FDC8",X"FDCE",X"FF8F",X"FF3A",X"FE06",X"FDC3",X"FD04",X"FDB2",X"FE9D",X"FE73",X"FCAB",X"F8E5",X"F52B",X"F2B6",X"F14E",X"F1A3",X"F2CE",X"FA1B",X"03B7",X"0BA1",X"102C",X"0F6E",X"0B1B",X"0567",X"FF7E",X"FD41",X"FD4F",X"FEE6",X"06E0",X"0D4A",X"0E3E",X"0AEC",X"03F7",X"FEE4",X"FE04",X"FDFF",X"FF0D",X"FDF6",X"FCC4",X"FC25",X"FBB8",X"FD50",X"FE8F",X"FE19",X"FC4F",X"F823",X"F4AD",X"F319",X"F217",X"F22C",X"F3E7",X"FAF9",X"03E5",X"0B58",X"0F6D",X"0DF2",X"0A01",X"0500",X"FFD5",X"FE01",X"FDDB",X"FF39",X"05BC",X"0BA1",X"0D0B",X"09DE",X"03CF",X"FF5F",X"FE42",X"FE6B",X"FF6E",X"FE48",X"FCEF",X"FC33",X"FB9A",X"FC64",X"FDBA",X"FD3F",X"FB35",X"F775",X"F40A",X"F2C5",X"F205",X"F15C",X"F424",X"FB35",X"02D6",X"09B5",X"0D73",X"0C6C",X"08E8",X"04DF",X"00F5",X"FF55",X"FF54",X"0162",X"070A",X"0BCA",X"0C62",X"0940",X"0366",X"00A4",X"0066",X"FF8D",X"FF6C",X"FE21",X"FC91",X"FC87",X"FC8F",X"FD8B",X"FEAA",X"FD30",X"FAB8",X"F73C",X"F401",X"F2E4",X"F2B6",X"F2C1",X"F6BF",X"FD5C",X"03CA",X"0980",X"0BFB",X"0B5C",X"08CA",X"051B",X"023F",X"00BC",X"003A",X"0233",X"0759",X"0B48",X"0B70",X"07A6",X"02EB",X"00BE",X"0004",X"FFCA",X"FF73",X"FDE1",X"FCAA",X"FC78",X"FD02",X"FE39",X"FEDA",X"FD70",X"FAE1",X"F74B",X"F4E8",X"F438",X"F409",X"F471",X"F7E0",X"FE6C",X"054C",X"09D4",X"0B7B",X"0A2A",X"0783",X"0551",X"03CD",X"02AF",X"02BB",X"04A9",X"08A6",X"0B3E",X"0A4A",X"070D",X"0371",X"01EB",X"0106",X"FFF3",X"FEE4",X"FD2D",X"FC2A",X"FBD0",X"FC3C",X"FD7C",X"FD90",X"FC01",X"F975",X"F608",X"F41D",X"F3A4",X"F391",X"F478",X"F890",X"FEA6",X"05A6",X"0974",X"0A09",X"08FC",X"0636",X"0468",X"0386",X"02B7",X"038B",X"048E",X"0710",X"087C",X"06C3",X"04AA",X"023F",X"0092",X"FFD0",X"FDF4",X"FCC7",X"FBE4",X"FB4C",X"FBCA",X"FCA6",X"FD03",X"FC0C",X"FA20",X"F80E",X"F548",X"F426",X"F497",X"F47E",X"F615",X"FA95",X"0030",X"0611",X"0816",X"082A",X"077D",X"0600",X"055B",X"0558",X"0551",X"0619",X"0682",X"06E0",X"06E8",X"053E",X"040E",X"034F",X"01CF",X"0093",X"FF33",X"FDC6",X"FCC0",X"FBF1",X"FC1F",X"FC5E",X"FBE6",X"FB2B",X"F98F",X"F745",X"F5CB",X"F4AB",X"F46F",X"F572",X"F8CA",X"FDFB",X"035A",X"068C",X"07DC",X"07E1",X"0730",X"06A9",X"05F4",X"0596",X"0570",X"0612",X"06A8",X"069B",X"05C8",X"049D",X"0350",X"0207",X"0099",X"FF3D",X"FDC9",X"FCD7",X"FC19",X"FC2C",X"FC9F",X"FC75",X"FBF2",X"FAFB",X"F93A",X"F775",X"F626",X"F5DF",X"F636",X"F812",X"FC71",X"013E",X"057B",X"07C1",X"078D",X"06C8",X"05CF",X"05B4",X"0647",X"06CC",X"067B",X"0597",X"04CA",X"04B7",X"0483",X"0420",X"02D0",X"0147",X"FF73",X"FE38",X"FD8C",X"FD31",X"FD2E",X"FD52",X"FCC0",X"FBDF",X"FB45",X"FA53",X"F8D9",X"F6EB",X"F63B",X"F676",X"F839",X"FC2D",X"0089",X"03FE",X"0655",X"073B",X"0731",X"06AD",X"06AF",X"06BC",X"06C7",X"0637",X"0528",X"04A1",X"0468",X"044E",X"042C",X"02EE",X"015E",X"FF8A",X"FDEF",X"FD49",X"FCC7",X"FC52",X"FC54",X"FC27",X"FB9A",X"FADA",X"F9D4",X"F859",X"F704",X"F659",X"F654",X"F7C6",X"FAD8",X"FEDC",X"029B",X"04A5",X"0578",X"05CF",X"059C",X"0555",X"0564",X"05BD",X"057C",X"04AD",X"03EC",X"0379",X"0357",X"030C",X"0292",X"01AF",X"FFE2",X"FE72",X"FDCC",X"FD99",X"FD8D",X"FD61",X"FCC5",X"FC05",X"FB9F",X"FB4D",X"FA46",X"F92F",X"F7E4",X"F6F9",X"F751",X"F986",X"FD37",X"012E",X"03C5",X"056E",X"065E",X"065A",X"05F2",X"05E5",X"05BF",X"0551",X"0463",X"03EE",X"0394",X"038D",X"036F",X"02F4",X"01E1",X"0074",X"FEEA",X"FE22",X"FD93",X"FD27",X"FCBD",X"FC38",X"FBA0",X"FB97",X"FB53",X"FA97",X"F994",X"F8AA",X"F80F",X"F871",X"FA2B",X"FD0C",X"0074",X"02EF",X"04A5",X"05F9",X"0686",X"06D0",X"06EC",X"073C",X"0719",X"05F7",X"0488",X"03AA",X"0379",X"03B6",X"0351",X"029C",X"013E",X"FFA4",X"FE80",X"FDEC",X"FD8C",X"FD38",X"FCAD",X"FBFB",X"FB33",X"FAF3",X"FADD",X"FA2B",X"F913",X"F841",X"F809",X"F960",X"FCA3",X"FFF8",X"022D",X"03A0",X"049F",X"0517",X"05BA",X"0689",X"0733",X"0736",X"0646",X"0500",X"0404",X"0397",X"03B1",X"0388",X"029C",X"0174",X"0043",X"FF48",X"FECE",X"FE8B",X"FDE8",X"FD32",X"FC22",X"FB04",X"FA9B",X"FAB5",X"FA4E",X"F9A9",X"F90E",X"F88D",X"F936",X"FB40",X"FE12",X"0093",X"0268",X"0374",X"03F6",X"0494",X"0507",X"05BA",X"0653",X"0605",X"0527",X"0411",X"034A",X"02FD",X"02D0",X"0268",X"0174",X"002D",X"FF33",X"FEBB",X"FEB4",X"FE76",X"FDB5",X"FC85",X"FB5E",X"FAAC",X"FA8B",X"FA3C",X"F9E1",X"F99C",X"F922",X"F8F7",X"FA99",X"FD86",X"0044",X"01D5",X"02B8",X"0370",X"042D",X"050C",X"05D0",X"0645",X"0611",X"051E",X"03ED",X"02E1",X"02B1",X"02C8",X"028D",X"0196",X"002D",X"FF4F",X"FECB",X"FE79",X"FE45",X"FD98",X"FC9C",X"FB97",X"FB09",X"FAB4",X"FA79",X"FA6E",X"FA18",X"F97D",X"F982",X"FA51",X"FC70",X"FF0D",X"0126",X"0231",X"02EF",X"03A8",X"049C",X"0585",X"065A",X"06B3",X"0647",X"0554",X"0456",X"03B9",X"0362",X"02F3",X"0206",X"00B1",X"FFAB",X"FF2D",X"FEFC",X"FEDC",X"FEA6",X"FDFF",X"FCE1",X"FBEF",X"FB75",X"FB01",X"FAC3",X"FAC3",X"FAB9",X"FAA2",X"FAB7",X"FC0A",X"FDF5",X"FFB9",X"00E7",X"01CE",X"02B5",X"035F",X"0416",X"04E3",X"0553",X"0568",X"0535",X"04BA",X"03E6",X"031A",X"02E0",X"02C0",X"0226",X"0162",X"0082",X"0011",X"FFC1",X"FF70",X"FEEA",X"FE19",X"FD60",X"FCE0",X"FC8B",X"FC6D",X"FC79",X"FC2E",X"FBEA",X"FB85",X"FB81",X"FCA1",X"FE6E",X"001D",X"0137",X"01C7",X"02A9",X"0387",X"043E",X"050B",X"0586",X"054E",X"04A7",X"040B",X"036D",X"032B",X"02E6",X"026C",X"0157",X"0031",X"FF59",X"FEB5",X"FE7B",X"FE51",X"FDE6",X"FD2E",X"FC4D",X"FBD5",X"FBA5",X"FBB1",X"FBC0",X"FB87",X"FB2C",X"FB53",X"FBC4",X"FCC1",X"FE24",X"FFD3",X"00F5",X"01B4",X"0227",X"02E0",X"03DC",X"047A",X"04D8",X"0511",X"049D",X"040A",X"034E",X"02C6",X"0284",X"022F",X"019C",X"00C8",X"FFD3",X"FF03",X"FE7D",X"FE59",X"FDFA",X"FD64",X"FC8B",X"FC0C",X"FBC8",X"FBCB",X"FC18",X"FC4C",X"FC32",X"FC68",X"FCC2",X"FD4C",X"FE55",X"FF81",X"00AC",X"018F",X"0232",X"02A4",X"02EE",X"038D",X"0421",X"048F",X"0478",X"03EA",X"0327",X"0266",X"01BD",X"013B",X"009B",X"FFDF",X"FF1C",X"FE7F",X"FDCD",X"FD89",X"FD50",X"FCCA",X"FC67",X"FC02",X"FBC5",X"FB80",X"FB80",X"FB86",X"FBAD",X"FC12",X"FC99",X"FD1B",X"FDEE",X"FF26",X"008C",X"01C4",X"02C0",X"039D",X"0447",X"048B",X"04CA",X"04F5",X"050C",X"04C9",X"043E",X"039B",X"02ED",X"025F",X"0201",X"0152",X"009E",X"FFE1",X"FF2A",X"FEDF",X"FE68",X"FDDD",X"FD79",X"FD15",X"FCF6",X"FCB0",X"FC96",X"FC85",X"FCDC",X"FD30",X"FD6F",X"FDA4",X"FE3C",X"FF80",X"009D",X"0135",X"0205",X"02A6",X"0330",X"0377",X"03E1",X"0419",X"03E8",X"0382",X"02E4",X"0237",X"0190",X"011B",X"00C9",X"0064",X"FFD5",X"FF4A",X"FEBE",X"FE49",X"FDF4",X"FDBC",X"FD88",X"FD50",X"FD42",X"FD0D",X"FCEF",X"FD0A",X"FD54",X"FD9F",X"FDF7",X"FE4D",X"FEBF",X"FFB9",X"0085",X"0137",X"01DE",X"02A3",X"0301",X"0303",X"033B",X"037A",X"038C",X"0382",X"0318",X"027A",X"01C5",X"0112",X"009E",X"0063",X"000A",X"FF9B",X"FF09",X"FE74",X"FDE6",X"FD59",X"FCFA",X"FCF4",X"FCDE",X"FCD2",X"FCAF",X"FCB2",X"FD04",X"FD16",X"FD5B",X"FDC9",X"FE52",X"FEF9",X"FF55",X"0012",X"00C8",X"01CA",X"025E",X"0234",X"023C",X"024D",X"02F2",X"031A",X"02C3",X"0281",X"020A",X"01EB",X"0113",X"0064",X"FF9C",X"FF4C",X"FF4B",X"FF24",X"FE8F",X"FE02",X"FDAD",X"FD2D",X"FCEF",X"FD05",X"FCEE",X"FD1B",X"FD95",X"FDE0",X"FDC2",X"FE03",X"FEA3",X"FF44",X"FF65",X"0006",X"004D",X"00C5",X"018B",X"021D",X"0247",X"021B",X"0225",X"024F",X"0267",X"0279",X"022B",X"0200",X"01C9",X"014B",X"00CD",X"0056",X"0009",X"FFAA",X"FF77",X"FF4C",X"FEEE",X"FE66",X"FE5B",X"FE20",X"FDFB",X"FDE6",X"FDFC",X"FE08",X"FE3D",X"FE78",X"FECA",X"FF77",X"0025",X"0086",X"00F5",X"0181",X"024D",X"02A0",X"031F",X"0369",X"0335",X"0303",X"02E0",X"0276",X"01E3",X"0148",X"00E8",X"00ED",X"0134",X"0111",X"00A6",X"003A",X"FFC1",X"FF0C",X"FEBE",X"FEC9",X"FE9D",X"FE53",X"FE11",X"FDFE",X"FE14",X"FE28",X"FDFB",X"FE30",X"FE7E",X"FEC7",X"FF0F",X"FF3B",X"FFB9",X"0014",X"0057",X"00A4",X"0117",X"01A9",X"01E6",X"01F9",X"01EF",X"01D1",X"01CB",X"0194",X"015E",X"012F",X"00E6",X"00F0",X"00B2",X"004D",X"0017",X"FF90",X"FF29",X"FEC2",X"FE59",X"FE04",X"FDD3",X"FDF5",X"FE00",X"FE0B",X"FE33",X"FE58",X"FE8C",X"FEC5",X"FF43",X"FF89",X"FFF1",X"0040",X"0093",X"00D6",X"00EC",X"0100",X"0100",X"0111",X"00F6",X"00FF",X"0124",X"00F6",X"007D",X"003A",X"0038",X"003F",X"0012",X"001C",X"FFE8",X"FF79",X"FF0C",X"FEC7",X"FE90",X"FE48",X"FE30",X"FE47",X"FE53",X"FE40",X"FE21",X"FE28",X"FE06",X"FDFF",X"FE68",X"FECB",X"FF0C",X"FF7B",X"FFC4",X"FFD2",X"FFF1",X"0022",X"0066",X"009B",X"009C",X"00A2",X"00A7",X"0066",X"004E",X"0043",X"0031",X"003D",X"0032",X"0011",X"000A",X"FFD6",X"FFAA",X"FFA1",X"FF94",X"FF6A",X"FF42",X"FF4B",X"FF3F",X"FF50",X"FF42",X"FF82",X"FF9C",X"FF9B",X"FFBE",X"FFED",X"0021",X"0021",X"0016",X"0050",X"009A",X"00D8",X"0103",X"0159",X"0181",X"0199",X"019D",X"016D",X"0162",X"016E",X"0160",X"0138",X"010D",X"00E8",X"00E2",X"00BA",X"0095",X"0055",X"0046",X"0035",X"001F",X"FFFA",X"FFC3",X"FFC7",X"FFD0",X"FFCE",X"FFD9",X"FFCE",X"FFBE",X"FF72",X"FF5C",X"FF7E",X"FF97",X"FFE1",X"0027",X"0066",X"0067",X"004F",X"0049",X"0034",X"0047",X"005A",X"006C",X"0071",X"0071",X"0072",X"0077",X"0051",X"000B",X"0013",X"0019",X"FFFF",X"FFDE",X"FF7D",X"FF41",X"FF3F",X"FF0B",X"FEDF",X"FECD",X"FF03",X"FF39",X"FF52",X"FF5E",X"FF47",X"FF1B",X"FF19",X"FF1A",X"FF44",X"FF8E",X"FF7A",X"FF98",X"FFD2",X"FFFE",X"0011",X"0059",X"0089",X"00A1",X"00A6",X"0070",X"0035",X"004B",X"0053",X"004D",X"005A",X"0042",X"0054",X"0058",X"0035",X"FFF5",X"FFAB",X"FF8D",X"FF64",X"FF35",X"FF27",X"FF08",X"FED5",X"FEF0",X"FF1D",X"FF4D",X"FF4B",X"FF94",X"FFD2",X"FFC6",X"FFC5",X"FFFD",X"0003",X"0012",X"004A",X"0064",X"0066",X"0084",X"007A",X"0068",X"005F",X"0070",X"0044",X"FFFC",X"0016",X"002E",X"FFF6",X"FFB7",X"FF88",X"FF92",X"FFAE",X"FFC5",X"FFC4",X"FFE4",X"FFCF",X"FFA7",X"FF7D",X"FF76",X"FF8E",X"FF66",X"FF74",X"FF91",X"FFA6",X"FF9E",X"FFBF",X"FFFD",X"002C",X"0031",X"0003",X"0008",X"0024",X"0034",X"004B",X"0041",X"0045",X"003C",X"0065",X"00A6",X"00BA",X"00AA",X"00A7",X"00A5",X"00A2",X"0088",X"004B",X"002A",X"0024",X"0015",X"0015",X"0036",X"0061",X"0030",X"001B",X"0020",X"FFF5",X"FFE8",X"FFFB",X"FFFC",X"0044",X"005E",X"005A",X"004A",X"0068",X"0088",X"00A2",X"00A7",X"0091",X"0074",X"002C",X"0009",X"002F",X"0043",X"0048",X"0016",X"0031",X"003B",X"0024",X"0012",X"FFF6",X"FFE0",X"FFE0",X"FF9E",X"FF70",X"FF76",X"FF85",X"FF65",X"FF6F",X"FF63",X"FF6A",X"FFAB",X"FFEA",X"FFD3",X"FFBA",X"FFCB",X"FFE8",X"FFFF",X"000A",X"FFFC",X"000E",X"000B",X"0035",X"006F",X"0090",X"007D",X"004B",X"003D",X"004F",X"0029",X"001E",X"0017",X"0012",X"0019",X"005C",X"0051",X"0022",X"0022",X"0009",X"FFF1",X"FFF4",X"FFED",X"FFBB",X"FFA1",X"FF84",X"FF64",X"FF38",X"FF3C",X"FF07",X"FEFF",X"FF34",X"FF48",X"FF5B",X"FF99",X"FFB9",X"0002",X"0026",X"0050",X"0049",X"004A",X"FFE8",X"FF7F",X"FF6C",X"FF84",X"FF8C",X"FF9A",X"FF3D",X"FF25",X"FF1D",X"FF42",X"FF33",X"FF0E",X"FF0E",X"FF0F",X"FF06",X"FEF5",X"FEBF",X"FEBF",X"FEC7",X"FEB4",X"FEDA",X"FF32",X"FF71",X"FF85",X"FF7A",X"FF7A",X"FF8F",X"FFB1",X"FFC7",X"FFF9",X"0016",X"0036",X"007B",X"00AD",X"009F",X"009C",X"00B2",X"00B3",X"0093",X"006A",X"006F",X"0072",X"0082",X"00AA",X"008E",X"007B",X"009B",X"00DA",X"00EB",X"00E9",X"00D3",X"0099",X"0062",X"0052",X"004D",X"0036",X"000F",X"0034",X"003C",X"0046",X"005B",X"005C",X"006F",X"0097",X"00CA",X"00E7",X"00DE",X"00B3",X"0083",X"009B",X"0095",X"0081",X"007C",X"0065",X"0058",X"006B",X"0055",X"0028",X"0001",X"FFB5",X"FF6D",X"FF76",X"FF7D",X"FF6F",X"FF9C",X"FFE2",X"FFED",X"FFEB",X"FFEA",X"FFF0",X"FFEC",X"0006",X"002F",X"0027",X"0025",X"0012",X"0011",X"002D",X"0029",X"0014",X"0019",X"0011",X"0057",X"006C",X"006F",X"0066",X"003F",X"000D",X"FFE2",X"FFB5",X"FFCA",X"FFDC",X"0000",X"0010",X"000A",X"0009",X"001B",X"0012",X"FFF2",X"FFED",X"FFB9",X"FFA1",X"FF9C",X"FFAA",X"FFA4",X"FF96",X"FF74",X"FF81",X"FF91",X"FF97",X"FF9F",X"FF8B",X"FF7E",X"FF93",X"FF7C",X"FF56",X"FF68",X"FFAE",X"FFC9",X"FFBB",X"FFA5",X"FFA1",X"FFC4",X"FFBF",X"FF91",X"FF5A",X"FF7F",X"FFC0",X"FFF3",X"FFED",X"FFC5",X"FFB3",X"FFC3",X"FFBE",X"FF93",X"FFB9",X"FFDE",X"FFF0",X"FFE9",X"FFCF",X"FFC4",X"FFCA",X"FFAD",X"FFAC",X"FFF2",X"FFF4",X"FFE0",X"FFE5",X"FFE7",X"FFBB",X"FF96",X"FFA8",X"FFB1",X"FFBC",X"FFA0",X"FF84",X"FF97",X"FFA3",X"FFAB",X"FFA8",X"FFBA",X"FFC1",X"FFBE",X"FFE1",X"FFFD",X"001B",X"001F",X"0041",X"0057",X"002C",X"001F",X"0023",X"0040",X"0078",X"0097",X"009F",X"00C6",X"00C1",X"00BA",X"00A2",X"0090",X"00B3",X"00B2",X"008C",X"004E",X"0057",X"00A7",X"00AC",X"0095",X"003F",X"0012",X"FFF0",X"FFEE",X"000B",X"001F",X"0019",X"FFEB",X"FFC7",X"FFB7",X"FF83",X"FFA1",X"FFF9",X"0017",X"0036",X"0022",X"FFFD",X"FFF1",X"FFA3",X"FF81",X"FF8A",X"FFB1",X"FFC0",X"FFF7",X"0004",X"FFEF",X"FFD0",X"FFAA",X"FF8C",X"FFAE",X"FFD1",X"0007",X"0010",X"001E",X"001D",X"FFD2",X"FFD0",X"000F",X"0039",X"002F",X"002C",X"002F",X"0001",X"0005",X"0001",X"FFF0",X"FFFE",X"0016",X"0068",X"0096",X"009E",X"0086",X"0090",X"0077",X"0068",X"006B",X"0058",X"0043",X"004C",X"003A",X"003D",X"0035",X"003B",X"003C",X"0034",X"0048",X"0018",X"FFCF",X"FFE1",X"0009",X"001A",X"FFF4",X"FFB8",X"FFBA",X"FFB0",X"FF93",X"FFA9",X"FFCA",X"FFBC",X"FFA0",X"FF87",X"FF73",X"FFC0",X"FFC1",X"FFC4",X"FFB5",X"FFAF",X"FFAE",X"FFC2",X"FFC8",X"FFBB",X"FFA6",X"FF90",X"FFA8",X"FFA9",X"FFC1",X"FF9B");
begin
 
   
 process(resetN, CLK)
	 type noteArrd is array (0 to 12) of integer;
	 variable dataTmp : noteArrd;
 begin
	if (resetN='0') then
		dataTmp := (others  => 0);
	elsif(rising_edge(CLK)) then
		dataTmp := (others  => 0);
		for i in 0 to 12 loop
			if conv_integer(addrArr(i)) > 0 then
				dataTmp(i) := conv_integer(sound0(conv_integer(addrArr(i))));
			end if;
		end loop;
	end if;
	Q <= conv_std_logic_vector(dataTmp(0) + dataTmp(1) + dataTmp(2) + dataTmp(3) + dataTmp(4) + dataTmp(5) + dataTmp(6) + dataTmp(7) + dataTmp(8) + dataTmp(9) + dataTmp(10) + dataTmp(11) + dataTmp(12), 16);
end process;
	 

		   
end arch;