--------------------------------------
-- SinTable.vhd
-- Written by Gadi and Eran Tuchman.
-- All rights reserved, Copyright 2009
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all ;

entity errtable is
port(
  CLK     					: in std_logic;
  resetN 					: in std_logic;
  ADDR    					: in std_logic_vector(14 downto 0);
  Q       					: out std_logic_vector(15 downto 0)
);
end errtable;

architecture arch of errtable is
constant array_size 			: integer := 2286 ;

type table_type is array(0 to array_size - 1) of std_logic_vector(15 downto 0);
signal err_table				: table_type;
signal Q_tmp       			:  std_logic_vector(15 downto 0) ;



begin
 
   
process(resetN, CLK)
	constant err_table : table_type := (X"F2F0",X"0A41",X"1000",X"F7AA",X"EAD1",X"EE2F",X"FFCD",X"1D31",X"0D1B",X"F686",X"EF7F",X"F418",X"0765",X"0692",X"0CA4",X"F6E8",X"05E7",X"023D",X"E044",X"FC32",X"05D1",X"106D",X"09DF",X"036A",X"03D7",X"1E7C",X"F977",X"E2FD",X"01E9",X"F8E4",X"FA28",X"FEB8",X"FF39",X"ECE3",X"F36B",X"00A8",X"0A25",X"18B5",X"0FD8",X"EFE7",X"E625",X"FB5D",X"FD54",X"1AB4",X"01FE",X"FEF1",X"0FCA",X"FAEE",X"F83F",X"0434",X"0C89",X"F932",X"0ADE",X"EF0E",X"F064",X"FEFD",X"095C",X"004F",X"ED12",X"0C16",X"1042",X"1FB8",X"F242",X"EC73",X"0E09",X"0075",X"F51F",X"F9BE",X"FF22",X"F6F7",X"18EE",X"F9B8",X"0592",X"1E8E",X"0D26",X"EF8E",X"F00D",X"021D",X"0A1E",X"1787",X"FD60",X"F90E",X"0434",X"02E3",X"06AE",X"0980",X"0C88",X"FBF1",X"0B3B",X"E7F3",X"E733",X"09FB",X"0AFE",X"0AAB",X"0F88",X"0919",X"0E24",X"0C88",X"E410",X"F05F",X"05DC",X"F883",X"FFA1",X"03CA",X"0FEC",X"0438",X"FD61",X"0007",X"0A34",X"1A2B",X"0725",X"EFF1",X"F5B3",X"FDE2",X"12CD",X"1143",X"F8DE",X"0614",X"107B",X"F13E",X"FED9",X"0AD3",X"0DEF",X"0EB4",X"F9AD",X"EB54",X"EBF9",X"0876",X"1464",X"02F2",X"02FF",X"1A14",X"1BE2",X"0944",X"EB5D",X"F905",X"00E5",X"EDDF",X"FEC5",X"0051",X"02F6",X"1543",X"09A7",X"0041",X"056C",X"12A2",X"0A67",X"F930",X"F0A3",X"0341",X"0AE1",X"0B08",X"0584",X"0103",X"034F",X"FD27",X"0394",X"03B3",X"056D",X"0CD5",X"F765",X"F0B3",X"ED51",X"FD1D",X"09FD",X"0F21",X"0D42",X"11CE",X"08CC",X"0269",X"F455",X"FD7C",X"F7D2",X"F23E",X"FDC3",X"068D",X"0477",X"00DD",X"03AF",X"039A",X"0A46",X"09CA",X"FB8A",X"F3D7",X"EF36",X"0287",X"0E16",X"06D2",X"047F",X"0D44",X"0324",X"F48F",X"0277",X"02A9",X"052D",X"123E",X"0311",X"F19F",X"F1FF",X"041C",X"09BF",X"06E1",X"0BA7",X"0A15",X"121F",X"FF2F",X"EE39",X"F331",X"F305",X"FBAA",X"0B57",X"058A",X"0222",X"0C07",X"01E2",X"F9FD",X"FC3B",X"FE15",X"03AB",X"F9F7",X"EE70",X"F25E",X"0E47",X"0EBD",X"FF60",X"FA84",X"F0C4",X"FCDE",X"117C",X"FFA4",X"F65A",X"FF40",X"F948",X"F69C",X"F601",X"FA4E",X"0F76",X"0973",X"0636",X"0155",X"087C",X"FB7A",X"F844",X"F8F8",X"E961",X"F52E",X"071D",X"0A12",X"069A",X"07DC",X"0503",X"06EF",X"07D8",X"FC88",X"FF47",X"EF8E",X"FE1B",X"00D0",X"0874",X"0292",X"0292",X"00DC",X"F7F1",X"0131",X"05D6",X"00D8",X"01B2",X"08EF",X"F968",X"F58A",X"FAD1",X"FC86",X"09E2",X"FBF8",X"007E",X"0563",X"123E",X"039C",X"F23A",X"EE33",X"F142",X"FA71",X"026F",X"055F",X"0615",X"08DE",X"FD1C",X"FACC",X"FEE4",X"FF52",X"0A49",X"FF5F",X"FD5B",X"F830",X"05A6",X"031C",X"00A9",X"FF51",X"F887",X"02D5",X"FBEE",X"FE16",X"FAAE",X"FCE9",X"FAFE",X"EF57",X"F9D7",X"FC68",X"0AFF",X"02A9",X"0558",X"037B",X"FF46",X"FDA2",X"F4E7",X"F2DD",X"EBCE",X"F14A",X"FC81",X"05F1",X"118A",X"001D",X"F9C2",X"FB55",X"004E",X"FB36",X"F871",X"F94C",X"FE93",X"FF29",X"0801",X"0D5B",X"078D",X"0621",X"FCA8",X"FA26",X"F517",X"021F",X"0D03",X"FE50",X"F55B",X"EF03",X"01CE",X"016D",X"0B74",X"020B",X"08F2",X"0FBD",X"07B5",X"00EB",X"F172",X"F81E",X"F3A0",X"F9CD",X"F91D",X"07D0",X"1729",X"02B9",X"F935",X"F0DD",X"FD4C",X"FDBC",X"0470",X"F9DC",X"F287",X"F6AD",X"02BC",X"001F",X"FDDA",X"051C",X"04F7",X"05EF",X"F2B8",X"F691",X"02EF",X"FD78",X"F592",X"EFF4",X"FCE9",X"FE72",X"0D74",X"00D8",X"FCF3",X"FD20",X"FEAB",X"F9F1",X"F141",X"F793",X"F8D3",X"018A",X"F804",X"FD39",X"0E53",X"0499",X"FD32",X"F69D",X"F9D4",X"F96B",X"033C",X"FD11",X"F3C8",X"FB3C",X"09FB",X"0053",X"FB81",X"FF8C",X"0612",X"00F5",X"F37F",X"F8F1",X"04E4",X"FE6D",X"EF31",X"F428",X"03E3",X"0578",X"0ACE",X"FF63",X"F8E2",X"FC79",X"04AD",X"FCC1",X"F475",X"EDEE",X"FA80",X"FA21",X"F71F",X"01FC",X"0DA4",X"07D4",X"F896",X"F999",X"F707",X"FEFB",X"04A0",X"F885",X"EEDC",X"FAFD",X"0B3D",X"01DE",X"FB4A",X"F8F9",X"0433",X"FFBF",X"F28F",X"F7DF",X"FEBB",X"FAFE",X"F2FA",X"FA99",X"0325",X"08B6",X"0A36",X"01F5",X"F800",X"FFA2",X"0055",X"FF50",X"FAA1",X"EFD7",X"F5D9",X"FB05",X"FD90",X"022F",X"0B9F",X"045D",X"FF3F",X"FDAA",X"F94F",X"02DA",X"05FB",X"FB50",X"F40B",X"FCE5",X"042A",X"00EF",X"054A",X"0449",X"057F",X"FF71",X"F461",X"FB02",X"FEA0",X"F26B",X"F358",X"FB9D",X"0310",X"067F",X"0A79",X"FC72",X"F62A",X"0063",X"FF63",X"04F4",X"F536",X"F3AD",X"F2D6",X"FA7C",X"00D0",X"0219",X"0925",X"FA83",X"F87E",X"F4F5",X"F4E0",X"034A",X"0033",X"F279",X"F4D8",X"0342",X"FFE1",X"0579",X"FFF3",X"FA68",X"FA7A",X"F8F5",X"F951",X"0442",X"0215",X"EBEB",X"F64F",X"FD21",X"09DB",X"0634",X"FF82",X"F804",X"FBBC",X"00E8",X"FCE3",X"0AB1",X"F83B",X"FDCA",X"FC35",X"FAB3",X"FF10",X"010D",X"0ECF",X"FE4E",X"0393",X"F811",X"FA0C",X"FFDE",X"F6BD",X"F82E",X"F97D",X"04BF",X"FEC9",X"0256",X"02D7",X"FF61",X"01C0",X"FB04",X"F83E",X"F8CC",X"F849",X"F0E0",X"FF7D",X"00AD",X"FDAD",X"030B",X"080F",X"FD84",X"FE56",X"004C",X"FE0B",X"0AA7",X"005F",X"F5AA",X"F32E",X"F452",X"FA83",X"02BD",X"08B8",X"FD46",X"0557",X"FFF6",X"F9B0",X"FB1F",X"F8D4",X"FCD4",X"FEFD",X"F7D4",X"FB4A",X"02E9",X"0AA6",X"FFA4",X"FBAB",X"F6D4",X"FE30",X"08BF",X"FD5C",X"F16B",X"FAB7",X"0780",X"04D8",X"05E6",X"004E",X"FF7A",X"005D",X"FFDA",X"FA54",X"FD12",X"FCE1",X"F6EB",X"FD21",X"F8A1",X"FB9E",X"080B",X"0584",X"FE14",X"FB6C",X"FC1A",X"FCE7",X"0188",X"FA58",X"FAF4",X"0366",X"FEF8",X"FD87",X"02FF",X"0634",X"FCD0",X"FCFA",X"F92B",X"FA9B",X"00FE",X"F909",X"F46F",X"FAE9",X"FDA2",X"016C",X"0898",X"0337",X"00A5",X"015D",X"F956",X"FB52",X"0031",X"0671",X"FBAA",X"0000",X"F72E",X"F834",X"028A",X"F9CC",X"F9E2",X"FBC5",X"F74A",X"F97A",X"FD39",X"F904",X"FA94",X"06D1",X"FC79",X"FA9E",X"00BD",X"0606",X"041F",X"FA4E",X"F214",X"F6E3",X"045C",X"FC59",X"F2CB",X"FABF",X"00C2",X"0892",X"0352",X"0096",X"FAF4",X"00DE",X"FD1B",X"F42E",X"FB4E",X"0020",X"00B9",X"0465",X"F919",X"F87B",X"034D",X"033C",X"01DE",X"FDC6",X"FC5F",X"078A",X"048A",X"FF09",X"F7F6",X"0640",X"FFA8",X"FFEE",X"FE36",X"0108",X"077E",X"06FF",X"FFD3",X"FBE1",X"0123",X"FCF6",X"FE21",X"FFE1",X"FB20",X"081E",X"0910",X"0563",X"FB9E",X"FBC3",X"F9A5",X"F9E1",X"FB59",X"FDBF",X"06F5",X"0A2C",X"0310",X"FD8D",X"FFB4",X"01BE",X"0637",X"FF6D",X"F756",X"029F",X"04E0",X"0357",X"0070",X"04AF",X"FF6E",X"019E",X"0038",X"FBBC",X"0488",X"012A",X"FEBD",X"F91E",X"FF54",X"0504",X"0726",X"05F7",X"FE78",X"06CF",X"06E7",X"033F",X"FE5C",X"0009",X"00A6",X"FFB2",X"FEA4",X"FDD1",X"06C6",X"0712",X"00BC",X"FB29",X"FEAF",X"0472",X"0430",X"FD67",X"F59C",X"FFC2",X"01D6",X"0268",X"FA20",X"024F",X"0360",X"00B4",X"0220",X"F9A4",X"01D9",X"0211",X"FCCA",X"F693",X"FA33",X"0552",X"02D8",X"FE84",X"F683",X"00B7",X"046A",X"0589",X"01C3",X"FB91",X"FB68",X"FA79",X"FD0B",X"F9A0",X"FFFE",X"03F1",X"FB0F",X"F4C5",X"F82E",X"012B",X"0470",X"FF7F",X"F92C",X"FFFB",X"01D4",X"03CA",X"01E9",X"FE5D",X"FE8A",X"FB8E",X"FF1C",X"F6AB",X"FC58",X"0109",X"FF5A",X"FDB0",X"FD49",X"036A",X"FFF2",X"FD46",X"F810",X"FC87",X"FFC0",X"0705",X"0ACE",X"02EC",X"00E9",X"00FC",X"018C",X"FCC0",X"FEFA",X"03CB",X"FA77",X"F9E6",X"FD56",X"04DF",X"FD26",X"FAE4",X"FA4D",X"FD71",X"0200",X"0127",X"031E",X"FD84",X"FE05",X"FF25",X"FF77",X"FD86",X"FD0E",X"029C",X"FC5C",X"FC76",X"FDD5",X"0691",X"0173",X"FD48",X"F988",X"F655",X"FE35",X"005C",X"05B0",X"FED5",X"FD1D",X"FFFA",X"FF94",X"FCE2",X"FE02",X"065A",X"FC60",X"FBD2",X"FC17",X"00AE",X"0266",X"03AF",X"0220",X"FFCF",X"0626",X"034B",X"0534",X"00A8",X"FEF2",X"00FA",X"04BA",X"FE21",X"FD44",X"0706",X"FFF8",X"FF16",X"0149",X"0291",X"0263",X"FE14",X"F981",X"F34D",X"FF09",X"0379",X"04D3",X"FEFE",X"F6D5",X"FE06",X"0174",X"FD2D",X"F8C4",X"FEF6",X"F9C2",X"FA8C",X"01EF",X"FC71",X"02AA",X"05C2",X"009B",X"FDEB",X"009F",X"0021",X"0320",X"FF7C",X"F935",X"FBB3",X"FED1",X"FFA7",X"FE91",X"02E4",X"FF73",X"0037",X"043D",X"FEA2",X"00D0",X"FF48",X"F947",X"F7DB",X"FA76",X"0037",X"0798",X"061E",X"00E0",X"01EC",X"00D6",X"FCE0",X"FF0C",X"023B",X"FE7A",X"FDED",X"FEC3",X"FD75",X"01BD",X"FF48",X"FCE1",X"0263",X"02DD",X"01CA",X"00C6",X"FD8B",X"F9CF",X"FD6C",X"FD5F",X"FA54",X"FEFF",X"01C2",X"0115",X"FF06",X"FEFA",X"FD2A",X"03A3",X"0223",X"FA9B",X"FE81",X"FFE9",X"042F",X"067B",X"0266",X"00DC",X"0439",X"01CF",X"FB6B",X"FCA7",X"FD0C",X"FD10",X"0029",X"FEC4",X"FD04",X"00CA",X"02BE",X"00C2",X"033C",X"FF6A",X"FF4D",X"00F9",X"FE36",X"FB71",X"FF13",X"FFED",X"FED6",X"FF69",X"0114",X"0251",X"02E1",X"0190",X"FE8D",X"FD2C",X"FB20",X"F92D",X"FF22",X"FE0F",X"0079",X"01C0",X"0204",X"008E",X"012D",X"020B",X"0035",X"0294",X"FFAD",X"FFD8",X"009E",X"003C",X"0202",X"FFC1",X"FEFE",X"FD02",X"0290",X"011B",X"01FA",X"00FE",X"FF32",X"FE49",X"FF3A",X"FE3D",X"FE51",X"016A",X"04B6",X"045E",X"02F8",X"FF34",X"FF8D",X"FF6B",X"FA47",X"FA17",X"FD78",X"FE30",X"0029",X"FFD9",X"FEF4",X"FFED",X"044A",X"0006",X"FB09",X"F8C7",X"F9E4",X"FEA0",X"FDEA",X"FD0A",X"FDFE",X"FDF5",X"FE23",X"FE77",X"0011",X"FC5B",X"FF42",X"0070",X"FE4F",X"FE12",X"FE87",X"FEFF",X"FF96",X"FE3E",X"FE1B",X"008E",X"03F5",X"0166",X"01D4",X"FE61",X"FCDD",X"0010",X"FF21",X"FEF3",X"0020",X"03B8",X"040A",X"02E9",X"0107",X"FCF1",X"FC8A",X"FA68",X"FECE",X"0206",X"013B",X"0214",X"00B9",X"0020",X"FEA2",X"023C",X"01BC",X"FEC0",X"FF40",X"0050",X"0317",X"01A6",X"FDDA",X"FBB8",X"FE04",X"014D",X"02D0",X"031A",X"0090",X"FEDB",X"FE23",X"FC12",X"FC16",X"FE5F",X"FFA9",X"005D",X"0134",X"03EC",X"0487",X"0508",X"02A0",X"FE05",X"FC39",X"FB3E",X"FE48",X"FF30",X"FF33",X"FEF1",X"FF0B",X"FFBE",X"001E",X"01F1",X"0039",X"FE31",X"FEEF",X"0102",X"01F2",X"FFBF",X"FC77",X"FC6A",X"FF01",X"0162",X"0237",X"02AA",X"0248",X"FF4B",X"FCD0",X"FB52",X"FFA1",X"0217",X"0207",X"0109",X"0236",X"0486",X"0528",X"05E2",X"0235",X"0110",X"FE69",X"FE3F",X"00EA",X"005C",X"0220",X"0146",X"004E",X"FF52",X"00D6",X"01A7",X"FFC2",X"FEDC",X"FE25",X"0217",X"0462",X"00A9",X"FB68",X"FC9C",X"FF8B",X"0229",X"04BC",X"025F",X"00C2",X"FE9A",X"FACB",X"FA76",X"FE04",X"016C",X"0282",X"01D6",X"012D",X"0212",X"033A",X"00E4",X"FDEA",X"FD20",X"FC09",X"FF40",X"0004",X"0018",X"00C9",X"00CC",X"FFAE",X"FF29",X"01CC",X"0048",X"FEC2",X"FAB6",X"FBAB",X"0141",X"035D",X"FF71",X"FC22",X"FEFB",X"01C5",X"054E",X"061A",X"040B",X"0150",X"FE7D",X"FBDF",X"FE01",X"00FF",X"038C",X"0454",X"0036",X"0000",X"035D",X"06BC",X"0264",X"FF10",X"FC7A",X"FC84",X"FFDD",X"FDE9",X"FF30",X"FFAF",X"FFBA",X"FFB0",X"0212",X"03FC",X"027E",X"01EF",X"FC19",X"FCBE",X"0188",X"0203",X"FECF",X"FC45",X"FC83",X"0014",X"03E1",X"02DE",X"00C6",X"FFA0",X"FBDB",X"FBA8",X"FCB0",X"FC64",X"FEF4",X"007B",X"FD6A",X"FDBA",X"FF3E",X"0098",X"FE55",X"FB39",X"F812",X"FC16",X"0029",X"FE85",X"FF10",X"FE4B",X"FDE7",X"FFD0",X"00AD",X"00D9",X"FFF9",X"FF6C",X"FB7E",X"FDF2",X"0179",X"0157",X"FFEC",X"FC33",X"FB2A",X"FE6C",X"0343",X"0304",X"FFA3",X"FC65",X"F8F5",X"FABD",X"FC8B",X"FD32",X"001A",X"0166",X"FF43",X"0036",X"01BA",X"00C7",X"002C",X"FD6D",X"FA5E",X"FCF0",X"007F",X"FF2C",X"0050",X"FFD8",X"FEF7",X"016A",X"0163",X"FF62",X"FF8B",X"FEFC",X"FCCB",X"FF96",X"0150",X"002C",X"0031",X"FDBB",X"FE06",X"014C",X"03DC",X"02E9",X"0194",X"FDC4",X"FC73",X"FE61",X"FCAE",X"FD21",X"01DC",X"0404",X"037D",X"0364",X"039C",X"0444",X"0429",X"FF68",X"FD98",X"011C",X"033A",X"0090",X"FE6B",X"FC52",X"FDC4",X"01B3",X"023B",X"0021",X"00BF",X"FF1B",X"FDD8",X"FF59",X"FEBF",X"00B2",X"022A",X"009B",X"FEFF",X"0120",X"0506",X"04D3",X"0265",X"FDB8",X"FE57",X"0102",X"010F",X"FFC0",X"00FA",X"01BD",X"0139",X"0174",X"0049",X"01F9",X"02CE",X"00DC",X"FEA0",X"0061",X"02FE",X"02A3",X"0109",X"FD79",X"FEEF",X"019F",X"0109",X"FFCE",X"FF27",X"FF4C",X"FF53",X"00D3",X"FEF9",X"008F",X"00C4",X"FEF4",X"FE9D",X"0093",X"0400",X"0330",X"0014",X"FBDF",X"FB7F",X"FDDC",X"FD01",X"FEC1",X"FFC8",X"012A",X"004D",X"FFB3",X"FEB0",X"FEBD",X"FE03",X"FB0B",X"FB95",X"FEB6",X"00FE",X"008E",X"FE2B",X"FF3A",X"01A9",X"0381",X"00C1",X"FFC5",X"FE8D",X"FDC7",X"FDCE",X"FE43",X"FDF8",X"00D0",X"01F1",X"FED4",X"FE1C",X"010C",X"0443",X"01DA",X"FD32",X"FC4C",X"FE39",X"FF84",X"FDDB",X"FE2A",X"FEC2",X"007D",X"00CB",X"002A",X"FE72",X"FFAB",X"00DF",X"FD1F",X"FDC0",X"FF55",X"0091",X"0023",X"FE6A",X"FE83",X"FFE7",X"01CF",X"00E7",X"008B",X"FFC3",X"FEA5",X"003F",X"FF90",X"FDC6",X"FFB2",X"0069",X"FE65",X"FF2C",X"0136",X"020A",X"00F3",X"FEE2",X"FCE9",X"FE61",X"FE08",X"FDB4",X"012D",X"0086",X"00E6",X"019A",X"00C5",X"FED7",X"FFF6",X"0155",X"FFB5",X"0219",X"01A7",X"0108",X"0053",X"FF13",X"FF7C",X"FFC2",X"FEBF",X"FED8",X"FFFD",X"FE38",X"FD04",X"FFC2",X"FF8B",X"FE4D",X"00C9",X"0161",X"0068",X"013A",X"021E",X"02C4",X"011C",X"0038",X"FEC4",X"FFF9",X"FECB",X"FF40",X"016E",X"0112",X"00FA",X"01AB",X"FF5C",X"FD0C",X"FEB6",X"FF4D",X"FE62",X"FF7A",X"FF3A",X"FF2A",X"FFBC",X"FEEC",X"FF0D",X"000C",X"FEFD",X"FECA",X"FF33",X"FD15",X"FCF8",X"FFEE",X"FE24",X"FC27",X"FDF6",X"FEB1",X"FF5E",X"0101",X"00B0",X"009A",X"0051",X"FD71",X"FD75",X"FCFA",X"FC2F",X"FDDE",X"FFEA",X"FF15",X"FE8A",X"0019",X"FF42",X"FE69",X"FFEA",X"0014",X"00DC",X"0212",X"0080",X"FF9C",X"0099",X"00E8",X"026E",X"0143",X"FFBE",X"00FC",X"02BD",X"0111",X"00BB",X"01B8",X"0132",X"0073",X"006C",X"FF69",X"FFD8",X"018B",X"00FD",X"0074",X"001B",X"FFC2",X"0161",X"FFEB",X"FD9C",X"FED4",X"0138",X"009A",X"00A6",X"0020",X"FEDC",X"FFBC",X"FFEC",X"FF6A",X"0104",X"018B",X"0073",X"000E",X"006A",X"0044",X"00C8",X"0025",X"FEFF",X"00F8",X"00C7",X"FF3E",X"FFAE",X"0026",X"FF87",X"0031",X"0011",X"FEF0",X"FFD6",X"006E",X"FFC4",X"FFE0",X"0032",X"FF2F",X"00C9",X"FECC",X"FDA3",X"FF62",X"00EE",X"003B",X"0017",X"002E",X"FF44",X"0012",X"FF4C",X"FEEF",X"0138",X"011C",X"FF57",X"FF4A",X"013A",X"019E",X"026E",X"FF51",X"FF1F",X"0087",X"0062",X"FEF0",X"FF96",X"FFC1",X"FF04",X"008C",X"FEE1",X"FF19",X"0128",X"01FB",X"018B",X"005D",X"FFD7",X"FF4C",X"014C",X"FEBD",X"FD70",X"FE7F",X"0061",X"0118",X"0016",X"FE11",X"FD12",X"FF0C",X"FE83",X"FEF9",X"0019",X"FF82",X"FDFE",X"FCE5",X"FE0F",X"FE3D",X"FFB3",X"FDAC",X"FDBF",X"FE41",X"FEAF",X"FF13",X"FFA0",X"FF45",X"FDCB",X"FF32",X"FEB8",X"FF55",X"FFFA",X"FFFF",X"FFDB",X"FEA2",X"FFB2",X"FF7C",X"014A",X"FFBD",X"FE8E",X"FEC7",X"FF88",X"00CE",X"FFEF",X"FEBD",X"FDAE",X"FF74",X"001D",X"0161",X"0291",X"0102",X"FED1",X"FE18",X"0038",X"00A5",X"00E7",X"FFDD",X"FFC5",X"FFE3",X"FFEA",X"FFF7",X"0003",X"FFBD",X"FF80",X"00B2",X"FFE4",X"0073",X"01D5",X"0158",X"000E",X"FF03",X"FFE1",X"0049",X"012C",X"FFB6",X"FE87",X"FF73",X"012D",X"01BE",X"0087",X"FEED",X"FE5F",X"FF02",X"FF95",X"0023",X"0120",X"0075",X"FE66",X"FDCC",X"FF1D",X"00A7",X"00E6",X"FFDA",X"FF1F",X"FEBD",X"FFA0",X"0085",X"0013",X"FEFF",X"FEC7",X"FF26",X"FF9F",X"FFCD",X"0138",X"011E",X"006B",X"FFB0",X"004F",X"0111",X"00D4",X"FFA7",X"FED8",X"FF69",X"00CF",X"0191",X"00B6",X"FFC0",X"0051",X"0095",X"0105",X"016B",X"01CF",X"00D6",X"FF61",X"FF22",X"0013",X"0210",X"0234",X"00C9",X"FFDC",X"FFEA",X"014D",X"0168",X"0094",X"FEEA",X"FF83",X"FFAF",X"FFB8",X"FFBA",X"00B7",X"00B3",X"0005",X"FF65",X"FF28",X"0103",X"0115",X"FF7A",X"FE53",X"FEBF",X"0031",X"00E2",X"FFCC",X"FD94",X"FE5E",X"FF32",X"0007",X"FFCB",X"0016",X"FF84",X"FEDA",X"FED6",X"FF08",X"00C0",X"010C",X"FFE4",X"FEA2",X"FE4C",X"FFBF",X"0089",X"001E",X"FE7D",X"FF84",X"0042",X"00F6",X"00D2",X"0109",X"0072",X"FF7F",X"FF31",X"FF20",X"008D",X"FFE5",X"FF16",X"FEF7",X"FF68",X"010C",X"016A",X"0068",X"FE74",X"FE9C",X"FEF1",X"FFD1",X"0078",X"0050",X"FF46",X"FEC6",X"FF52",X"0046",X"0199",X"015B",X"FFFD",X"FF46",X"FF2A",X"FFD9",X"0000",X"FF80",X"FE61",X"FF2E",X"FF65",X"004E",X"00E3",X"00FE",X"003E",X"FF87",X"FF2E",X"FF42",X"007D",X"FFEC",X"FEF7",X"FED8",X"FF1C",X"007D",X"0056",X"FF64",X"FE5E",X"FED3",X"FFCC",X"00BD",X"00A5",X"FFFC",X"FE9F",X"FE4D",X"FECD",X"FFBE",X"011C",X"00AE",X"FF87",X"FEE6",X"FF1C",X"FFF5",X"0022",X"FFBA",X"FEFD",X"FF51",X"FF4A",X"0027",X"0047",X"FFE5",X"FF2E",X"FED6",X"FF16",X"FFC5",X"009B",X"00B6",X"0024",X"0008",X"0032",X"00C3",X"00D1",X"FFB5",X"FEBB",X"FEDC",X"FF9A",X"00A2",X"0094",X"FF9F",X"FEB6",X"FF24",X"FFD4",X"00EF",X"0137",X"00C5",X"FFBF",X"FF07",X"FEEB",X"FF8A",X"0058",X"0028",X"FFB4",X"FF62",X"FF81",X"00D2",X"0121",X"0058",X"FF2B",X"FEA7",X"FEBE",X"FF73",X"FF93",X"FFE1",X"FFA0",X"FF63",X"FFF4",X"00BB",X"00B4",X"FFEE",X"FF59",X"FF30",X"FF91",X"0068",X"0076",X"FFA3",X"FF38",X"FF54",X"FFD6",X"00FA",X"00F1",X"00C0",X"FFE4",X"FF62",X"FF7C",X"0038",X"009A",X"006E",X"0024",X"FF9B",X"0031",X"011C",X"0104",X"0051",X"FFC6",X"FFA4",X"FFB9",X"0026",X"0043",X"0046",X"FFE6",X"FFAA",X"FFDE",X"009F",X"00AF",X"0015",X"FF58",X"FF16",X"0017",X"00D8",X"00AB",X"FFD9",X"FF8B",X"FF95",X"0005",X"0036",X"0006",X"0015",X"FFA9",X"FF46",X"FF42",X"0013",X"00A0",X"0091",X"001B",X"FF66",X"FFF6",X"00E8",X"00CA",X"FFFC",X"FF55",X"FF3A",X"FF99",X"000C",X"0000",X"000E",X"FFF8",X"FFE1",X"0009",X"0054",X"0050",X"FFC8",X"FF2B",X"FEF1",X"FF82",X"0044",X"0029",X"FFC3",X"FF99",X"FF5F",X"FFDF",X"0085",X"0089",X"004D",X"FFC7",X"FF8C",X"FFA6",X"FFE8",X"0019",X"FFEF",X"0006",X"003B",X"00BA",X"0115",X"00F8",X"0070",X"FFE5",X"FF98",X"FFA0",X"FFEB",X"002E",X"0046",X"0011",X"FFDC",X"0036",X"00CE",X"009E",X"FFD5",X"FF50",X"FF71",X"0016",X"0036",X"FFED",X"FFBA",X"FFB7",X"FFA0",X"FFE4",X"002A",X"0028",X"0003",X"FF9B",X"FF4F",X"FF74",X"FFF4",X"0022",X"FFCE",X"FF95",X"FF73",X"FFC9",X"0032",X"0049",X"FFE5",X"FF97",X"FFA5",X"0021",X"002F",X"0020",X"FFF8",X"FFB5",X"FFA5",X"FFB5",X"FFE7",X"FFC7",X"FF7F",X"FF40",X"FF4A",X"FFD0",X"002F",X"003B",X"FFEF",X"FFCC",X"FF93",X"FFC8",X"FFFF",X"0004",X"FFD1",X"FF8A",X"FF95",X"0000",X"004E",X"004A",X"001D",X"FFD7",X"FFB7",X"FFB1",X"FFE6",X"002D",X"0026",X"FFEE",X"FFB6",X"000E",X"0026",X"0062",X"0041",X"FFFC",X"0000",X"0047",X"0066",X"001B",X"FFE0",X"FFA6",X"FFCE",X"0015",X"0019",X"001A",X"000C",X"001B",X"0018",X"0036",X"0049",X"007B",X"005A",X"0003",X"FFC0",X"0007",X"003C",X"002B",X"FFEA",X"FFA4",X"FFB7",X"FFEC",X"001E",X"0025",X"FFE6",X"FFCC",X"FFCF",X"FFD2",X"FFC7",X"FFE3",X"FFE0",X"FFE5",X"FFEF",X"0008",X"0023",X"0003",X"FFD8",X"FFB6",X"FFB1",X"FFD2",X"FFF4",X"FFFA",X"FFD4",X"FFB4",X"FFAB",X"FFE5",X"0015",X"0045",X"0011",X"FFE4",X"FFD9",X"0016",X"0032",X"0015",X"0010",X"FFF0",X"FFFD",X"0026",X"0038",X"004C",X"0029",X"000C",X"FFDE",X"FFEA",X"000B",X"0041",X"0033",X"FFE3",X"FFEC",X"0002",X"0021",X"000A",X"FFDE",X"FFE1",X"FFEC",X"0013",X"000C",X"FFFB",X"0008",X"000C",X"0002",X"FFFE",X"0013",X"002A",X"000C",X"FFD7",X"FFD3",X"000F",X"0030",X"001E",X"FFF5",X"FFD8",X"FFE3",X"FFEF",X"0002",X"000D",X"FFF9",X"FFF3",X"FFD8",X"FFCD",X"FFD6",X"FFF6",X"0000",X"FFF2",X"FFEC",X"FFEC",X"FFF2",X"FFDC",X"FFC2",X"FFC8",X"FFD3",X"FFF4",X"FFF9",X"FFF8",X"FFF4",X"0009",X"0008",X"0003",X"0014",X"001A",X"0005",X"FFED",X"FFF5",X"0008",X"0012",X"0001",X"FFF3",X"FFED",X"FFED",X"FFF6",X"0003",X"0004",X"0007",X"0006",X"FFF2",X"FFE4",X"FFEF",X"0005",X"0006",X"0004",X"0007",X"000C",X"0014",X"000A",X"0004",X"FFFD",X"0003",X"0005",X"0006",X"FFFD",X"FFFA",X"FFFB",X"FFEF",X"FFEB",X"FFF7",X"0000",X"FFFA",X"FFF5",X"FFF9",X"0000",X"0000",X"FFF8",X"FFEE",X"FFEC",X"FFED",X"FFF0",X"FFF2",X"FFF2",X"FFF9",X"FFF9",X"FFF8",X"FFF7",X"FFFB",X"FFFF",X"FFFF",X"0000",X"FFFE",X"0001",X"0000",X"FFFF");
begin
	if (resetN='0') then
		Q_tmp <= ( others => '0');
	elsif(rising_edge(CLK)) then
	--      if (ENA='1') then
		Q_tmp <= err_table(conv_integer(ADDR));
	--      end if;
	end if;
end process;

Q <= Q_tmp; 

		   
end arch;