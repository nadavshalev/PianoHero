--------------------------------------
-- SinTable.vhd
-- Written by Gadi and Eran Tuchman.
-- All rights reserved, Copyright 2009
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all ;

entity metronomTable is
port(
  CLK     					: in std_logic;
  resetN 					: in std_logic;
  ADDR    					: in std_logic_vector(9 downto 0);
  Q       					: out std_logic_vector(15 downto 0)
);
end metronomTable;

architecture arch of metronomTable is
constant array_size 			: integer := 601 ;

type table_type is array(0 to array_size - 1) of std_logic_vector(15 downto 0);
signal Q_tmp       			:  std_logic_vector(15 downto 0) ;



begin
 
   
process(resetN, CLK)
	constant metronom_table : table_type := (X"0024",X"001F",X"0019",X"0011",X"0004",X"FFFB",X"FFF7",X"FFF0",X"FFEF",X"FFF4",X"FFFA",X"FFFB",X"FFFF",X"0013",X"0018",X"001A",X"0023",X"0034",X"0030",X"0036",X"0048",X"0045",X"0040",X"003D",X"004C",X"005E",X"0059",X"0051",X"004F",X"0060",X"0074",X"0065",X"0062",X"006C",X"0059",X"004D",X"004D",X"004C",X"003C",X"0034",X"0034",X"0034",X"0033",X"0043",X"006E",X"0059",X"003D",X"0069",X"0092",X"0060",X"0071",X"004A",X"0079",X"0057",X"003F",X"0067",X"0084",X"006B",X"0094",X"0054",X"007C",X"009F",X"0056",X"0057",X"0092",X"0093",X"0065",X"00B7",X"007B",X"008C",X"006E",X"007E",X"00B4",X"00D7",X"0070",X"00B8",X"0116",X"00E0",X"00AA",X"0075",X"00F7",X"01A6",X"0161",X"00FF",X"0107",X"00F0",X"01DC",X"01A7",X"0153",X"0200",X"026D",X"02D2",X"028D",X"02C6",X"035E",X"0315",X"02A4",X"037E",X"0426",X"02EB",X"033A",X"03E7",X"0366",X"0271",X"0247",X"0221",X"01F8",X"00BD",X"0033",X"0037",X"0079",X"FF96",X"FF2A",X"FD2E",X"FDA5",X"FD58",X"FCEA",X"FC83",X"FB25",X"FBF7",X"FCF1",X"FB01",X"FA8C",X"FB36",X"FA8E",X"FB50",X"FA4A",X"F9F9",X"FB4A",X"FB85",X"FB2A",X"FAFB",X"FAF1",X"FC24",X"FD89",X"FC6D",X"FCDB",X"FD88",X"FD56",X"FEFE",X"FF3D",X"FE80",X"FEEF",X"FD76",X"F851",X"FBFE",X"FADD",X"F3CC",X"F3DC",X"F52B",X"FE08",X"0754",X"DE99",X"F10B",X"CCA2",X"F9D7",X"403F",X"3C21",X"F546",X"C706",X"3671",X"4414",X"18DB",X"DE75",X"C48F",X"C4FB",X"16AB",X"393F",X"261E",X"E3B6",X"CB7C",X"E117",X"FEB2",X"2E1F",X"0946",X"02CB",X"DCD3",X"EDBA",X"FD68",X"167F",X"0C0B",X"0515",X"FABD",X"01BC",X"F8EC",X"0104",X"0151",X"0EA4",X"08EC",X"084F",X"F9A0",X"FB0B",X"FDEE",X"0A29",X"0EC5",X"09B4",X"00BE",X"FBA5",X"FEE1",X"0743",X"0B7D",X"092E",X"0398",X"0069",X"FE4C",X"03BB",X"0688",X"0762",X"06E7",X"02CA",X"017F",X"FE58",X"0567",X"06E5",X"052D",X"0764",X"033C",X"FEEE",X"0317",X"06EA",X"0754",X"0608",X"02E8",X"00D8",X"FEED",X"0417",X"07D8",X"0532",X"0038",X"FFDB",X"0093",X"034C",X"02BB",X"041B",X"02B2",X"FE78",X"0022",X"01F6",X"0331",X"0359",X"017D",X"FF73",X"0060",X"02CF",X"026C",X"029A",X"01A4",X"0084",X"01A5",X"00DC",X"00DB",X"01BE",X"0071",X"010B",X"009B",X"0131",X"FFB9",X"FF99",X"FE52",X"0177",X"0231",X"0162",X"0097",X"FF56",X"FF0B",X"0083",X"0196",X"0101",X"0131",X"0019",X"FF69",X"FFC8",X"FED2",X"FF19",X"00E5",X"023C",X"01C0",X"0018",X"FCB7",X"FDDD",X"01CC",X"0235",X"041F",X"002F",X"FCEE",X"FE9D",X"FFDE",X"02BB",X"010A",X"0074",X"FDEE",X"FD8A",X"FFE3",X"0174",X"0273",X"FF8A",X"FDE2",X"FD45",X"FFAE",X"0198",X"009B",X"FF6A",X"FE5A",X"FEE7",X"FF88",X"00E7",X"FFB5",X"FF8C",X"FF02",X"FF6B",X"FF9C",X"0082",X"FF53",X"FEDF",X"FFA7",X"FF88",X"002D",X"FDEA",X"FCD5",X"FF22",X"FF73",X"FF72",X"FE73",X"FCD4",X"FFAF",X"0058",X"0007",X"FD1F",X"FCE9",X"FE40",X"FE18",X"00DD",X"FF32",X"FDAA",X"FEA9",X"FEB4",X"FF59",X"FF11",X"FDC3",X"FDCD",X"FF43",X"FE73",X"FEF8",X"FFCD",X"FB16",X"0027",X"FF11",X"0014",X"FEDB",X"FEA8",X"FEDB",X"024E",X"FD0A",X"FC80",X"FF06",X"FD36",X"0335",X"FE0A",X"FE12",X"FC40",X"FE77",X"0179",X"00A7",X"FDEC",X"FEB1",X"FC44",X"0065",X"010E",X"FEE0",X"013B",X"0090",X"FD64",X"FE5A",X"FECC",X"00E0",X"01CE",X"FFBF",X"FF76",X"FF60",X"FC0D",X"0206",X"00A3",X"FEA0",X"00D3",X"FCE9",X"00D0",X"FE41",X"01C3",X"002A",X"0003",X"00BE",X"FDAC",X"FFA5",X"FE87",X"042F",X"02B1",X"00CA",X"FE2D",X"FE93",X"FF65",X"02FC",X"0021",X"FD53",X"FA07",X"FD92",X"051B",X"0688",X"036D",X"FE0F",X"FB7A",X"FC79",X"0182",X"00A7",X"FD25",X"00F0",X"01C8",X"0203",X"0206",X"FD6F",X"FE93",X"0048",X"02E2",X"0061",X"FE6B",X"F75F",X"FF93",X"015E",X"047A",X"041D",X"FD9B",X"FD48",X"00F8",X"018D",X"0209",X"FDC8",X"FEF3",X"FF47",X"0178",X"023B",X"FE67",X"FDD4",X"00C5",X"01F3",X"0266",X"FF71",X"FC4F",X"FC58",X"0027",X"0252",X"0383",X"00DF",X"FDAC",X"FE32",X"FFD4",X"01EA",X"01A9",X"010E",X"FE29",X"FCDD",X"FD45",X"FFA0",X"0084",X"020B",X"017B",X"00AE",X"FFE8",X"FEE6",X"FFA5",X"FF83",X"FF93",X"00A3",X"0158",X"FF8A",X"FE39",X"FEB7",X"0045",X"FF64",X"02B4",X"FE53",X"FFAB",X"FE2F",X"FEBB",X"0147",X"FECB",X"008E",X"FEE1",X"0143",X"0092",X"00A0",X"FEFD",X"FDAB",X"FFD0",X"011C",X"016C",X"00FF",X"FE67",X"FC4D",X"00D4",X"FFC2",X"037D",X"FFBD",X"FF74",X"FF71",X"FE8E",X"0059",X"01C0",X"016F",X"FF3A",X"FDC9",X"FE32",X"FF1B",X"0165",X"0165",X"00E5",X"FDFE",X"FE35",X"FCA7",X"00FF",X"0137",X"00AD",X"0086",X"FF4E",X"FEA1",X"FF24",X"FFBF",X"FF53",X"FFD4",X"00D7",X"0060",X"FEB8",X"FE61",X"01CC",X"FFBB",X"007E",X"FF01",X"FFAF",X"FF5F",X"0193",X"FDF1",X"FCFD",X"FC30",X"019D",X"0188",X"0123",X"FE6D",X"FD9A",X"FFCD",X"00B2",X"0153",X"0137",X"FDAF",X"FF1D",X"FFA0",X"FFDF",X"00AB",X"FFBD",X"FE6F",X"FF58",X"00DF",X"0106",X"FF6D",X"FF74",X"002A",X"FFC1",X"010B",X"FFC0",X"FF10",X"FF53",X"0037",X"00A6",X"00E6",X"006F",X"FFCA",X"FF63",X"005E",X"FF7C",X"0031",X"0067",X"FFCA",X"FF48",X"FEC5",X"FF6F",X"FFA1",X"0005",X"00B1",X"00DA",X"FF4B",X"0033",X"FFBF",X"FF44",X"000B",X"014E",X"012B",X"FFCC",X"FEEA",X"FF98",X"FF78",X"0136",X"00DE",X"FFDE",X"002D");
begin
	if (resetN='0') then
		Q_tmp <= ( others => '0');
	elsif(rising_edge(CLK)) then
		Q_tmp <= metronom_table(conv_integer(ADDR));
	end if;
end process;

Q <= Q_tmp; 

		   
end arch;