library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_signed.all ;
use ieee.std_logic_arith.all;
library work;
use work.pkg2.all;

package pkg2 is
  type Arr_type is array (0 to 12) of std_logic_vector(13 downto 0);
end package;

package body pkg2 is
end package body;


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_signed.all ;
use ieee.std_logic_arith.all;
library work;
use work.pkg2.all;

entity piano_effect is
port(
  CLK     					: in std_logic;
  resetN 					: in std_logic;
  addrArr    				: in Arr_type;
  Q       					: out std_logic_vector(15 downto 0)
);
end piano_effect;

architecture arch of piano_effect is
	constant array_size 			: integer := 8201 ;
	
	signal Q_tmp       			:  std_logic_vector(15 downto 0) ;
	
	type table_type is array(0 to array_size - 1) of std_logic_vector(15 downto 0);
	constant sound0 : table_type := (X"0008",X"FFF8",X"0006",X"FFFF",X"0000",X"0007",X"FFFF",X"FFF7",X"0007",X"0006",X"FFF4",X"FFF4",X"FFF8",X"FFFB",X"0000",X"FFF8",X"FFF7",X"FFF9",X"FFFE",X"FFFF",X"FFFF",X"0000",X"0004",X"FFFB",X"0008",X"FFFF",X"0004",X"FFFC",X"FFFD",X"0000",X"0008",X"0004",X"000A",X"0007",X"000F",X"0001",X"FFF5",X"0002",X"0002",X"FFFB",X"0000",X"0000",X"0005",X"0001",X"FFF4",X"0000",X"FFF4",X"FFF2",X"FFFD",X"FFF9",X"FFF7",X"0004",X"0005",X"0002",X"0004",X"FFFE",X"0006",X"0000",X"0007",X"0009",X"0001",X"0002",X"0005",X"0008",X"FFFE",X"FFF8",X"FFF7",X"0000",X"FFF7",X"FFFA",X"0004",X"0003",X"0001",X"FFFE",X"0006",X"FFFC",X"0002",X"000D",X"FFFC",X"0002",X"FFF9",X"0000",X"0000",X"FFFF",X"0005",X"0001",X"FFFF",X"FFF8",X"0000",X"FFFF",X"FFEE",X"FFF6",X"FFF2",X"0002",X"FFFF",X"FFFD",X"FFFB",X"0001",X"0008",X"0006",X"0005",X"0004",X"0000",X"FFF5",X"0007",X"0009",X"FFFB",X"0000",X"0008",X"0000",X"FFF9",X"0000",X"FFF7",X"0000",X"0000",X"FFFE",X"0000",X"FFF7",X"FFF8",X"FFFC",X"0001",X"FFFE",X"FFF6",X"FFFB",X"FFFB",X"FFFA",X"FFF8",X"FFF0",X"FFFC",X"0000",X"000B",X"000F",X"0004",X"0000",X"0001",X"FFFC",X"000E",X"FFF7",X"FFF9",X"0005",X"FFFB",X"0003",X"0001",X"FFF8",X"FFF8",X"FFF7",X"FFF9",X"FFF9",X"FFFA",X"0001",X"0000",X"0003",X"0000",X"FFFF",X"0000",X"0004",X"FFF8",X"0008",X"0005",X"FFF8",X"0004",X"FFFC",X"0004",X"FFFA",X"FFFA",X"0001",X"FFFE",X"0007",X"0000",X"0003",X"0000",X"0001",X"FFFE",X"FFF7",X"FFF0",X"0000",X"0007",X"0002",X"FFFB",X"0000",X"0008",X"0002",X"FFFC",X"FFFE",X"FFFD",X"0002",X"0003",X"0002",X"FFFB",X"0003",X"0001",X"0003",X"0000",X"000B",X"FFF8",X"FFF5",X"0004",X"000B",X"0006",X"0003",X"FFFB",X"FFF1",X"FFFF",X"0010",X"FFFE",X"0005",X"FFF8",X"FFF6",X"FFFE",X"0000",X"0008",X"FFFB",X"0004",X"0000",X"0001",X"FFFF",X"FFFA",X"0000",X"FFF5",X"FFFB",X"0001",X"FFF8",X"FFFD",X"FFFC",X"000F",X"FFFF",X"FFFF",X"0000",X"FFFD",X"0002",X"0000",X"0004",X"0000",X"FFFA",X"FFFD",X"FFFA",X"000B",X"0008",X"0007",X"000E",X"0000",X"FFF6",X"0000",X"0007",X"FFFE",X"0004",X"FFFB",X"FFFE",X"FFF7",X"FFF9",X"FFFE",X"0006",X"0007",X"FFFF",X"0000",X"FFF6",X"0000",X"FFFD",X"0003",X"0001",X"0008",X"0003",X"FFF9",X"000A",X"0009",X"000B",X"0007",X"0008",X"0003",X"FFF8",X"FFF8",X"FFF5",X"FFFE",X"0008",X"FFF6",X"0001",X"0001",X"FFF9",X"FFFB",X"FFFD",X"0000",X"0003",X"0000",X"0000",X"0002",X"0001",X"FFFF",X"0009",X"0005",X"FFFC",X"FFF9",X"FFF3",X"0001",X"FFFF",X"FFF6",X"FFED",X"FFF5",X"FFFD",X"0003",X"000E",X"FFFA",X"0007",X"FFFA",X"0000",X"0009",X"0000",X"0000",X"FFF3",X"FFFA",X"FFF1",X"0002",X"FFF6",X"FFFD",X"FFFE",X"FFFA",X"0002",X"0003",X"0005",X"FFFD",X"FFFE",X"FFFF",X"0000",X"0001",X"FFFB",X"FFFD",X"0001",X"0001",X"0004",X"FFF8",X"0000",X"0014",X"000B",X"000C",X"FFF9",X"FFFE",X"0004",X"FFFF",X"0000",X"0006",X"0005",X"0000",X"FFFA",X"FFFB",X"000C",X"0001",X"FFFD",X"0000",X"0006",X"000A",X"FFFF",X"FFFD",X"0004",X"0001",X"0008",X"0000",X"FFFB",X"FFF3",X"FFFF",X"FFF4",X"FFEF",X"0006",X"0000",X"0005",X"0006",X"FFFF",X"FFFE",X"0001",X"000B",X"0005",X"FFFF",X"0000",X"FFFE",X"FFF7",X"FFF8",X"FFFD",X"0003",X"0005",X"0005",X"0000",X"FFF7",X"FFF6",X"FFF4",X"0006",X"0000",X"0002",X"0003",X"FFFE",X"FFFD",X"FFF6",X"0001",X"0006",X"0004",X"FFFE",X"0000",X"FFFE",X"0004",X"0007",X"0001",X"FFFC",X"FFFF",X"0002",X"0004",X"FFF9",X"0005",X"0005",X"0000",X"0001",X"FFFD",X"FFFE",X"0000",X"0001",X"FFF6",X"FFFC",X"0007",X"FFFE",X"0000",X"000A",X"0002",X"0002",X"0000",X"0001",X"FFF8",X"FFFD",X"0007",X"FFF2",X"FFF7",X"FFF7",X"FFFB",X"FFFA",X"0001",X"0000",X"0002",X"0009",X"FFFC",X"0004",X"0007",X"0004",X"0009",X"FFFA",X"0003",X"FFF8",X"0001",X"0003",X"0004",X"0008",X"0000",X"000C",X"0004",X"FFFE",X"FFF9",X"FFFB",X"0000",X"0001",X"FFFC",X"0001",X"FFF9",X"FFF7",X"0004",X"0001",X"0000",X"0009",X"FFFD",X"FFF5",X"FFF9",X"FFF8",X"0002",X"0000",X"FFFE",X"000C",X"000A",X"0003",X"FFFE",X"FFFC",X"0000",X"0004",X"0003",X"0000",X"0002",X"FFFE",X"FFF2",X"FFFF",X"000B",X"0007",X"FFFE",X"FFFE",X"FFFF",X"0007",X"0004",X"0007",X"0001",X"FFF3",X"FFEF",X"FFFC",X"FFFB",X"FFFE",X"FFF5",X"0004",X"FFF3",X"0001",X"0007",X"0002",X"0008",X"000C",X"000C",X"0008",X"0009",X"000C",X"0002",X"FFF8",X"0000",X"0001",X"FFF8",X"FFF9",X"FFF1",X"FFF8",X"FFF8",X"FFFD",X"FFFC",X"0003",X"FFFD",X"FFF9",X"0005",X"0000",X"FFF4",X"FFF5",X"0003",X"000F",X"0007",X"000C",X"0005",X"0001",X"0006",X"FFFB",X"FFF9",X"0000",X"FFFB",X"0000",X"0003",X"000A",X"0000",X"FFF9",X"0001",X"0002",X"FFFC",X"FFFD",X"0001",X"0009",X"FFF4",X"FFEF",X"FFF7",X"0009",X"0006",X"0017",X"0001",X"FFFE",X"0007",X"FFFE",X"000C",X"0005",X"0003",X"0003",X"FFFA",X"FFF5",X"FFF1",X"000B",X"0001",X"FFF5",X"000D",X"0001",X"0008",X"FFFD",X"0006",X"FFF8",X"FFF0",X"FFED",X"FFFB",X"FFF2",X"0000",X"0002",X"0005",X"0009",X"0003",X"FFFC",X"0006",X"0007",X"FFFD",X"0009",X"000B",X"0007",X"FFF2",X"FFFE",X"FFF7",X"FFFB",X"FFFE",X"FFF9",X"FFFA",X"0009",X"FFFE",X"FFF4",X"0005",X"0007",X"0000",X"FFFE",X"000B",X"0009",X"FFF9",X"FFF4",X"0003",X"FFF3",X"FFEA",X"FFF4",X"FFFE",X"0007",X"0007",X"0012",X"000E",X"0003",X"FFF8",X"0010",X"000A",X"FFF8",X"FFFB",X"0008",X"FFF9",X"FFED",X"FFF9",X"FFF2",X"0009",X"FFFB",X"000C",X"0019",X"0004",X"0002",X"0000",X"FFF8",X"0000",X"0009",X"FFF9",X"0005",X"0010",X"0000",X"0003",X"0004",X"0006",X"FFEE",X"FFFD",X"0004",X"FFF6",X"FFF1",X"0002",X"0005",X"0000",X"FFF3",X"0004",X"0015",X"0005",X"0002",X"000B",X"0007",X"0000",X"FFFC",X"0004",X"0003",X"FFF0",X"FFFB",X"0004",X"FFF5",X"FFFB",X"FFFC",X"0005",X"0000",X"000E",X"0018",X"000C",X"000C",X"FFF6",X"FFFA",X"FFFD",X"FFF6",X"FFFE",X"0008",X"0002",X"FFFF",X"FFFD",X"FFFE",X"0003",X"FFFE",X"0004",X"0011",X"0011",X"0003",X"FFFD",X"FFFC",X"FFF8",X"FFF6",X"0001",X"000B",X"FFE8",X"FFF2",X"FFFD",X"FFE1",X"FFDB",X"FFEB",X"FFF4",X"FFE6",X"FFEE",X"0006",X"0002",X"FFFD",X"002B",X"0029",X"002C",X"003F",X"0041",X"004A",X"003A",X"0057",X"004A",X"004F",X"0036",X"FEFD",X"FEA2",X"FFB9",X"FFFC",X"0024",X"FF92",X"FEC2",X"0166",X"0395",X"0310",X"0312",X"010D",X"00E1",X"FE2D",X"FA0C",X"F3E5",X"F06A",X"F607",X"F896",X"00B6",X"0E2F",X"1832",X"1B6E",X"1848",X"0F7A",X"FB61",X"EC13",X"E59D",X"E7EE",X"F1A2",X"F7CC",X"FCB5",X"0231",X"0B70",X"0DD0",X"0A94",X"0CDD",X"0BC6",X"0370",X"023C",X"02E3",X"FAF3",X"F0C3",X"E59D",X"E361",X"EFA3",X"F7FE",X"FFA3",X"09DA",X"18B1",X"1FED",X"1A52",X"1AD4",X"1A28",X"0889",X"F2F5",X"EE3C",X"ECE0",X"EA51",X"E211",X"D6C0",X"E186",X"F48A",X"067B",X"16E1",X"253B",X"2B34",X"2025",X"0FBA",X"052A",X"FE05",X"F178",X"EB63",X"F14F",X"F8A7",X"FA73",X"EAB5",X"E00E",X"E5A6",X"F215",X"01D5",X"174D",X"2B1C",X"2FDB",X"27EA",X"1C1B",X"0D82",X"F6CE",X"E1DA",X"E040",X"E661",X"EDDE",X"E68F",X"DA87",X"E6E7",X"FD87",X"0C5C",X"19E6",X"2C54",X"35C1",X"2A3D",X"146A",X"FE54",X"ED1F",X"DBE2",X"D82E",X"E704",X"FC88",X"031C",X"F06F",X"E918",X"F853",X"0476",X"073D",X"0F47",X"1E0A",X"22C0",X"1C30",X"0E90",X"008D",X"F491",X"EE53",X"F3B1",X"FCA1",X"0077",X"EEEE",X"DCB6",X"E7D9",X"FD25",X"02F9",X"040F",X"0F03",X"18DE",X"19CA",X"14BF",X"0C75",X"03F3",X"F841",X"F4D0",X"F8C0",X"FF3B",X"F661",X"DDC5",X"D878",X"EEB3",X"0287",X"066A",X"0D8C",X"1AC6",X"1F84",X"1BAE",X"1302",X"0B20",X"FF5F",X"F6FC",X"F3CE",X"F6A1",X"F98D",X"E85B",X"D5C5",X"E21A",X"FE13",X"09DB",X"0AEA",X"1346",X"17F0",X"170C",X"11FC",X"0A48",X"FF95",X"F7AC",X"F85B",X"FD41",X"072F",X"01E0",X"E7AD",X"DD04",X"EE38",X"FCB5",X"FB03",X"FFFE",X"0BA3",X"12D3",X"1597",X"13B0",X"0C4C",X"0067",X"FB30",X"FAB9",X"033E",X"0C04",X"FD18",X"E400",X"E3B1",X"F54A",X"F9AE",X"F875",X"0100",X"09AB",X"1068",X"139D",X"1434",X"0CFD",X"04B2",X"FDD0",X"FC2B",X"0835",X"0881",X"EDDF",X"D937",X"E1A5",X"EE10",X"F048",X"FBEA",X"0BDF",X"1832",X"1D0D",X"1E1B",X"1963",X"0D71",X"0003",X"F1C5",X"F43E",X"0315",X"FC17",X"E5B2",X"E42A",X"F584",X"F956",X"F86C",X"FEEA",X"07AD",X"0E8A",X"11B4",X"135B",X"0DBB",X"0719",X"FDF0",X"F9A6",X"0922",X"1153",X"FBF4",X"E4DE",X"E79D",X"ED9A",X"EB35",X"F0C4",X"FD39",X"0B13",X"126F",X"17AB",X"1578",X"0EC6",X"066E",X"F9E5",X"FDE0",X"1058",X"0C88",X"F138",X"E4A0",X"EBDB",X"EC8F",X"ECEF",X"F3F1",X"01A7",X"0D75",X"15D0",X"192E",X"14B9",X"0ED3",X"0277",X"F995",X"069D",X"1196",X"FE2C",X"E245",X"DFD3",X"E4C0",X"E574",X"EADF",X"F912",X"0AF7",X"187F",X"224A",X"219D",X"1AFE",X"0F2E",X"FC92",X"FA23",X"0A06",X"09A8",X"EED9",X"DEDB",X"E2E3",X"E5D8",X"E7FE",X"EF28",X"FEDE",X"0C70",X"1803",X"1D6B",X"19DF",X"1459",X"0631",X"F99A",X"0390",X"1213",X"0536",X"EB7F",X"E5F1",X"E89E",X"EA53",X"EC9E",X"F5F3",X"01A6",X"0C62",X"1675",X"1730",X"1477",X"0D47",X"FD31",X"FAB4",X"0D08",X"1287",X"F9CE",X"E6A4",X"E3F6",X"E5B7",X"E7CE",X"EF73",X"FDA6",X"0A3E",X"1700",X"1D2E",X"1C05",X"19B1",X"0BCE",X"FB22",X"FFBB",X"0F1A",X"0439",X"EA35",X"DECB",X"DD80",X"DEF9",X"E389",X"F110",X"01C0",X"1325",X"2282",X"2578",X"239C",X"1AE3",X"05D6",X"F984",X"04D0",X"098A",X"F2FD",X"DF37",X"DAC9",X"DF08",X"E51A",X"F137",X"01BC",X"108E",X"1ED5",X"2323",X"1EC8",X"193E",X"089C",X"F2DF",X"F281",X"0461",X"00C9",X"EE01",X"E40C",X"E665",X"EBE4",X"F227",X"FCEF",X"078A",X"130F",X"1C03",X"1ACC",X"17C5",X"1010",X"FBAC",X"ECC4",X"FAA7",X"082F",X"FD98",X"ED62",X"E7A3",X"EA9E",X"EE52",X"F510",X"FE4B",X"08DE",X"15F2",X"1B29",X"193D",X"16EE",X"0A42",X"F32A",X"F0C3",X"0468",X"0803",X"F9A1",X"ED81",X"EC1A",X"ED86",X"EF6A",X"F500",X"FB8F",X"06CC",X"1226",X"14F2",X"16E9",X"156A",X"048F",X"F370",X"FE89",X"0D27",X"072F",X"F70A",X"EE39",X"EC89",X"EADC",X"ED50",X"F29A",X"FB9F",X"0A8A",X"13D3",X"1739",X"1A8E",X"1468",X"FD8C",X"F6B5",X"054C",X"0A1E",X"FCBC",X"EE3F",X"EA74",X"EA32",X"EC48",X"F207",X"F8CC",X"0554",X"11E7",X"1692",X"18A4",X"1A7B",X"0A59",X"F5E2",X"FB38",X"085C",X"049F",X"F426",X"EA1F",X"E8BD",X"E9CD",X"EF96",X"F5DC",X"FE50",X"0BFA",X"1537",X"17E2",X"1C5E",X"1810",X"00E2",X"F5C2",X"00E7",X"0826",X"FD95",X"EEA9",X"E98F",X"E97F",X"EC60",X"F158",X"F5D5",X"00E4",X"0DC1",X"142E",X"18CB",X"1EDC",X"1107",X"FAA7",X"FA6F",X"0770",X"0802",X"F92F",X"ED4B",X"E940",X"E827",X"EBA8",X"EF3D",X"F7B8",X"068B",X"12B1",X"1739",X"1F3D",X"1E8E",X"0772",X"F719",X"FDDA",X"07CD",X"0092",X"F166",X"E977",X"E71C",X"EA3C",X"EF46",X"F470",X"FFB4",X"0E4A",X"14CC",X"1933",X"2143",X"158E",X"FDB6",X"F74C",X"0297",X"066B",X"F9D4",X"ED84",X"E8B4",X"E912",X"ED34",X"EFC7",X"F5EC",X"03A6",X"100B",X"14BA",X"1EB7",X"212B",X"0D7B",X"FA68",X"FC93",X"06C8",X"036C",X"F5FC",X"ECE0",X"E899",X"E9EB",X"EBD4",X"EE90",X"F810",X"07EE",X"100D",X"1727",X"2202",X"1AA7",X"03AF",X"F8A8",X"019E",X"0863",X"FF58",X"F375",X"EC01",X"EB2C",X"EDC5",X"EFB5",X"F2BF",X"FE78",X"0A22",X"0E79",X"1973",X"1FC9",X"10F2",X"FCA2",X"FAFB",X"062E",X"066B",X"FB70",X"F106",X"EBF9",X"EC76",X"EE6A",X"EF1B",X"F523",X"0313",X"0A25",X"11D3",X"1F51",X"1E3B",X"09E6",X"FADC",X"FF84",X"06E6",X"0116",X"F5B2",X"ED07",X"EB25",X"ED0A",X"EEBF",X"F06B",X"FC22",X"07DB",X"0CC4",X"17EF",X"214D",X"15FA",X"FFE3",X"F8D4",X"02BA",X"063F",X"FEEE",X"F469",X"EE4E",X"ED6C",X"EF77",X"EF0C",X"F3BB",X"00B7",X"0761",X"0DBE",X"1B3E",X"1DFD",X"0C24",X"FA3D",X"FCE6",X"05A8",X"046A",X"FB0C",X"F220",X"EE76",X"F031",X"F16A",X"F0D3",X"FA51",X"0428",X"0719",X"1051",X"1CA2",X"1721",X"01CB",X"F8AF",X"008D",X"0699",X"02A4",X"F932",X"F227",X"F0AE",X"F2E3",X"F019",X"F1F8",X"FCC3",X"02A9",X"076C",X"159D",X"1D7E",X"0FB0",X"FD19",X"FCD7",X"05F5",X"0881",X"012A",X"F74E",X"F082",X"F07E",X"EF61",X"EC5D",X"F411",X"FEA5",X"02CB",X"0CDD",X"1C31",X"1C37",X"089B",X"FC6A",X"0119",X"0821",X"05DA",X"FC4C",X"F296",X"EF06",X"F079",X"ECC4",X"EDEE",X"F8EE",X"FFBC",X"04D3",X"135A",X"1F90",X"15A2",X"0286",X"FD9E",X"04CD",X"089C",X"02FE",X"F946",X"F11E",X"F15F",X"F04C",X"EC62",X"F251",X"FBDF",X"FFC5",X"0823",X"18A3",X"1CAE",X"0BE3",X"FD2D",X"FEFC",X"07B2",X"08CF",X"0211",X"F76E",X"F232",X"F1E0",X"ED01",X"EC77",X"F5C4",X"FC22",X"003E",X"0DAC",X"1D01",X"181F",X"05F9",X"FD9E",X"0398",X"0915",X"0673",X"FD33",X"F3E8",X"F28C",X"F068",X"EAF5",X"EF6F",X"F90E",X"FCBB",X"033A",X"1546",X"1ED0",X"1278",X"01EE",X"FFF3",X"073C",X"098C",X"0420",X"F864",X"F23E",X"F1DB",X"EC1B",X"E9C7",X"F250",X"F9D2",X"FC88",X"093B",X"1BC5",X"1C9D",X"0C19",X"0041",X"0322",X"0868",X"089B",X"FFFB",X"F5AE",X"F36F",X"F0D3",X"EA4F",X"ECE9",X"F6A1",X"FA68",X"FF09",X"10A1",X"1E27",X"1691",X"0584",X"0062",X"04CE",X"08C7",X"05AE",X"FAA9",X"F439",X"F3B4",X"EE3E",X"EA70",X"F159",X"F8B1",X"FA49",X"04FD",X"184E",X"1E5F",X"10E9",X"034D",X"0231",X"067E",X"0824",X"0050",X"F574",X"F31C",X"F0DA",X"EA6C",X"EBAE",X"F593",X"FA0F",X"FDD5",X"0E22",X"1E4A",X"1B31",X"0A67",X"0197",X"02EC",X"076C",X"0632",X"FBD4",X"F516",X"F3FC",X"EE82",X"E93F",X"EF06",X"F730",X"F906",X"01DC",X"14EA",X"1F34",X"1469",X"05E3",X"01A8",X"050C",X"08E1",X"0354",X"F947",X"F5F6",X"F34B",X"EBD3",X"EAFA",X"F3E0",X"F7E3",X"F9C4",X"070B",X"19A3",X"1B5F",X"0D8B",X"0307",X"01EF",X"06DC",X"07AE",X"FEA7",X"F74F",X"F597",X"F080",X"EA91",X"EF46",X"F720",X"F880",X"FE82",X"10C3",X"1E8D",X"1811",X"0978",X"011F",X"01F8",X"0657",X"023B",X"F902",X"F5A1",X"F461",X"EDF4",X"EBF7",X"F3E1",X"F88A",X"F9AA",X"0471",X"17C5",X"1D12",X"112A",X"041F",X"FF6A",X"041E",X"073E",X"00F2",X"FA50",X"F8EE",X"F43B",X"EC37",X"EE12",X"F4C5",X"F632",X"F8CC",X"0910",X"1991",X"17F1",X"0B72",X"019D",X"01DC",X"0827",X"0731",X"FF67",X"FB8C",X"F9E2",X"F1C1",X"ECAD",X"F13E",X"F573",X"F432",X"FBB6",X"0F09",X"1955",X"1354",X"0790",X"0118",X"04D9",X"090C",X"03F7",X"FCF1",X"FB4A",X"F6BA",X"EE11",X"ED9E",X"F3B4",X"F4FF",X"F543",X"0387",X"15F9",X"19BC",X"106D",X"049C",X"01D6",X"06E0",X"06DB",X"0009",X"FBEF",X"FA7B",X"F26C",X"EC0A",X"EF31",X"F440",X"F2D9",X"F85B",X"0B50",X"18F9",X"175B",X"0BE7",X"0318",X"0509",X"096B",X"05B7",X"FEA3",X"FD0C",X"F86A",X"EF3F",X"EC4D",X"F191",X"F317",X"F1B8",X"FDA6",X"10B4",X"18F7",X"12E4",X"0701",X"02AD",X"074B",X"0907",X"02CA",X"FEB1",X"FCDF",X"F588",X"EDAD",X"EED4",X"F3DD",X"F216",X"F4BB",X"0510",X"14B6",X"1750",X"0E10",X"0426",X"045F",X"092D",X"06C5",X"006C",X"FE7B",X"FA91",X"F17C",X"EC9B",X"F0CC",X"F2A1",X"F025",X"F947",X"0BC0",X"17C4",X"15EA",X"0B10",X"04CF",X"07D6",X"09E8",X"03EF",X"FF83",X"FD7E",X"F6C0",X"ED90",X"ECF1",X"F1F3",X"F02A",X"F176",X"FFFE",X"11A9",X"18FB",X"1273",X"07E0",X"0549",X"09A0",X"07A8",X"01CA",X"FF7C",X"FC6F",X"F396",X"ECE5",X"F06F",X"F23F",X"EF29",X"F554",X"066D",X"1518",X"16DC",X"0D4D",X"04BF",X"06B7",X"096B",X"04B1",X"0042",X"FEB4",X"F979",X"EFD6",X"EE4B",X"F32E",X"F1CE",X"F0F5",X"FC1B",X"0D78",X"1805",X"1494",X"0968",X"0489",X"07E1",X"0688",X"00EA",X"FE62",X"FCEF",X"F584",X"EE73",X"F18E",X"F40A",X"F0D1",X"F41B",X"0270",X"1294",X"17BA",X"0FCD",X"057D",X"054C",X"07E5",X"048C",X"00C5",X"0025",X"FCC3",X"F2F4",X"EFAC",X"F32F",X"F186",X"EF02",X"F696",X"077A",X"14BE",X"152E",X"0AE8",X"04FE",X"07C3",X"07AF",X"0365",X"00F6",X"0088",X"F968",X"F147",X"F282",X"F453",X"F0A5",X"F0B9",X"FC38",X"0C9A",X"1583",X"1059",X"0626",X"04E0",X"079A",X"059B",X"01B1",X"01A2",X"FF2B",X"F5BE",X"F163",X"F44F",X"F38F",X"F012",X"F440",X"02EA",X"11B6",X"1585",X"0C6C",X"0526",X"0644",X"06E7",X"035A",X"0130",X"01AE",X"FB98",X"F2F2",X"F293",X"F454",X"F142",X"EF59",X"F7F7",X"07EE",X"142C",X"1275",X"08F2",X"05E8",X"07AA",X"06C6",X"0313",X"0360",X"01E9",X"F8DF",X"F2EE",X"F3F3",X"F335",X"EE80",X"EFE5",X"FC12",X"0C69",X"13FC",X"0D90",X"0683",X"0686",X"087D",X"05AA",X"03CC",X"04E3",X"FF7D",X"F649",X"F388",X"F47B",X"F0FF",X"ED5C",X"F2C6",X"01D7",X"10E5",X"129D",X"0AC7",X"067A",X"0824",X"07B8",X"03E8",X"0427",X"034A",X"FAE1",X"F3DA",X"F3CB",X"F396",X"EF40",X"EEDF",X"F887",X"0966",X"1416",X"104E",X"088E",X"0689",X"07ED",X"0517",X"030F",X"049A",X"006E",X"F7C7",X"F401",X"F4CE",X"F21A",X"EE16",X"F0AE",X"FDAE",X"0DF3",X"128C",X"0C6B",X"06EA",X"07D1",X"07E3",X"04B8",X"0581",X"0578",X"FE59",X"F669",X"F4E1",X"F418",X"EF73",X"ECF1",X"F305",X"036E",X"1048",X"104D",X"095C",X"06DA",X"08B6",X"069A",X"04FB",X"06AE",X"03B6",X"FAF4",X"F58C",X"F51B",X"F23F",X"EDB0",X"ED49",X"F84B",X"0969",X"1211",X"0E76",X"0899",X"08BE",X"08A0",X"0536",X"0566",X"0605",X"0005",X"F7C2",X"F514",X"F44A",X"F08B",X"ECB5",X"F031",X"FF5A",X"0E60",X"11D4",X"0BA6",X"07B7",X"0894",X"062E",X"0442",X"060B",X"04C9",X"FCFD",X"F6E0",X"F5F4",X"F3AE",X"EF14",X"EC58",X"F4E7",X"0592",X"10E8",X"0FA2",X"0950",X"0856",X"07E6",X"04D0",X"04B3",X"0636",X"01CD",X"F9B8",X"F698",X"F595",X"F2B6",X"ED9B",X"EE98",X"FB77",X"0BA4",X"1241",X"0D1F",X"0857",X"081E",X"05B5",X"033D",X"04C7",X"04A5",X"FDBE",X"F80A",X"F692",X"F592",X"F185",X"ED2C",X"F2B3",X"020E",X"0FC9",X"1115",X"0AC5",X"087E",X"075C",X"040A",X"0363",X"0578",X"029C",X"FB50",X"F78C",X"F679",X"F48B",X"EECE",X"ED38",X"F735",X"07B0",X"1183",X"0E97",X"09F7",X"08FA",X"066D",X"036D",X"0479",X"055E",X"FF87",X"F9CA",X"F734",X"F68E",X"F2A5",X"ED13",X"EFAC",X"FCF4",X"0C95",X"10DE",X"0C35",X"0966",X"07B5",X"03FF",X"0262",X"0524",X"0379",X"FDCC",X"F9B0",X"F8AC",X"F753",X"F159",X"ED56",X"F384",X"02D1",X"0EA6",X"0E38",X"09FC",X"0847",X"05B3",X"0257",X"03C3",X"059E",X"0213",X"FCA9",X"F97A",X"F8FB",X"F539",X"EEA8",X"EDD4",X"F854",X"0863",X"0F61",X"0CC0",X"09FA",X"081B",X"044B",X"0250",X"04DC",X"0452",X"FF8A",X"FA9A",X"F93F",X"F840",X"F2A1",X"ED4B",X"F078",X"FE97",X"0C20",X"0E8A",X"0BAB",X"09CC",X"0752",X"0346",X"03F1",X"0577",X"02F1",X"FD90",X"F9BA",X"F961",X"F65D",X"EFE8",X"EC91",X"F44D",X"0413",X"0D67",X"0D54",X"0B05",X"096A",X"0525",X"02D9",X"04D4",X"0560",X"01E3",X"FC7F",X"FA82",X"F972",X"F468",X"EDA7",X"ED93",X"F9A0",X"080C",X"0D31",X"0BF0",X"0AB2",X"07EA",X"0387",X"0394",X"05A9",X"04F8",X"0008",X"FBAB",X"FAC5",X"F838",X"F1BA",X"EC31",X"F0D2",X"FF7A",X"0A7E",X"0C91",X"0B4D",X"0A2A",X"05B4",X"02F2",X"046A",X"05FD",X"03AA",X"FE24",X"FB7E",X"FA59",X"F610",X"EEF9",X"EC2E",X"F5EF",X"0465",X"0BF0",X"0C1C",X"0BB5",X"08CA",X"0422",X"035C",X"0545",X"05D2",X"0173",X"FCD1",X"FB5D",X"F957",X"F3C7",X"EC9A",X"EE59",X"FB02",X"079B",X"0BE2",X"0C2D",X"0B5F",X"06DB",X"0392",X"0402",X"063C",X"04B7",X"FF85",X"FC69",X"FB21",X"F7E2",X"F0AA",X"EB9A",X"F210",X"FFE3",X"0941",X"0BA0",X"0C71",X"0A10",X"059C",X"03BB",X"0531",X"066D",X"02B8",X"FE20",X"FC2C",X"FA79",X"F5A1",X"ED88",X"EC80",X"F6D5",X"042A",X"0A60",X"0C63",X"0C5F",X"0874",X"04B8",X"03F7",X"0614",X"0522",X"0040",X"FD0B",X"FBB2",X"F9AC",X"F29B",X"EC28",X"EF92",X"FC75",X"06F8",X"0B03",X"0CD1",X"0AE5",X"06CD",X"03DD",X"04B3",X"0638",X"0322",X"FF05",X"FCCB",X"FBFD",X"F7EC",X"EFB5",X"EBDF",X"F39B",X"008F",X"0801",X"0BAB",X"0C64",X"099F",X"0571",X"03BC",X"05DD",X"05A9",X"01AA",X"FE37",X"FCF5",X"FBAF",X"F538",X"ED5A",X"ED67",X"F890",X"036D",X"0948",X"0C70",X"0BDC",X"0826",X"042D",X"044B",X"0634",X"03EF",X"0021",X"FD65",X"FD18",X"FA03",X"F23E",X"EC0E",X"F0DE",X"FCC1",X"0577",X"0ADA",X"0CBC",X"0AD8",X"0665",X"0395",X"0575",X"05A0",X"02A7",X"FEC4",X"FD75",X"FCAF",X"F7BE",X"EF4D",X"EC9A",X"F54B",X"FFBF",X"076E",X"0BFF",X"0C80",X"0968",X"04D6",X"0463",X"05DD",X"04BC",X"00E6",X"FDFE",X"FDB6",X"FBC5",X"F4F1",X"ED20",X"EF68",X"F947",X"0296",X"093D",X"0C4E",X"0BAC",X"0744",X"03E8",X"04E9",X"0555",X"0319",X"FF48",X"FE0B",X"FDD6",X"FA67",X"F1C8",X"ED38",X"F342",X"FCF8",X"0555",X"0ABD",X"0C81",X"0A28",X"0503",X"03E6",X"0502",X"04A9",X"013E",X"FE82",X"FE5B",X"FDB1",X"F7ED",X"EF41",X"EF14",X"F6C5",X"FFD6",X"0748",X"0B38",X"0BDC",X"0777",X"03E8",X"0425",X"0521",X"0399",X"002C",X"FEE0",X"FEF4",X"FD0A",X"F4AC",X"EE9C",X"F1B3",X"F9C3",X"0251",X"083A",X"0B99",X"0A2A",X"0595",X"03F7",X"0506",X"0579",X"0289",X"FFD8",X"FF00",X"FF46",X"FA55",X"F16A",X"EEB9",X"F3E9",X"FCA5",X"0499",X"09F8",X"0C25",X"0884",X"04B5",X"042A",X"0574",X"0433",X"010A",X"FEB0",X"FEE0",X"FE17",X"F6C0",X"EFBB",X"F074",X"F72C",X"0001",X"06CB",X"0BDB",X"0B2A",X"06C0",X"0403",X"04AB",X"0552",X"0304",X"0036",X"FED6",X"FFC5",X"FC13",X"F382",X"EF56",X"F242",X"FA65",X"0239",X"08D4",X"0C2A",X"0980",X"056B",X"0420",X"056A",X"0480",X"01EE",X"FF2B",X"FF68",X"FF51",X"F8B2",X"F13F",X"EF8F",X"F4C8",X"FCE6",X"044A",X"0A9F",X"0B9C",X"082A",X"04D4",X"0534",X"0572",X"03C9",X"00B9",X"FF0E",X"0045",X"FD9A",X"F5A0",X"F005",X"F0B5",X"F7C6",X"FF69",X"0716",X"0B9A",X"0A6E",X"065D",X"048E",X"0525",X"04B2",X"0293",X"FFC1",X"0018",X"00CC",X"FB32",X"F3A3",X"EF8C",X"F2FB",X"F9EE",X"0184",X"08AA",X"0B1E",X"0894",X"0538",X"0501",X"055D",X"0497",X"01D1",X"FFEE",X"016C",X"FF44",X"F839",X"F133",X"EFF3",X"F517",X"FC16",X"0447",X"0A36",X"0AF1",X"075F",X"0560",X"0579",X"0563",X"039C",X"0067",X"0081",X"0151",X"FCE6",X"F565",X"EFFA",X"F18F",X"F6FE",X"FE98",X"0686",X"0B28",X"09BF",X"0683",X"059C",X"05DA",X"0553",X"0242",X"FFE1",X"0136",X"FFEF",X"FA34",X"F2AB",X"EFFE",X"F31B",X"F967",X"01BB",X"0925",X"0B85",X"089C",X"0648",X"05C6",X"05DE",X"0465",X"0096",X"0069",X"0138",X"FE4F",X"F740",X"F0E7",X"F08D",X"F4A8",X"FC05",X"0498",X"0AD9",X"0A9B",X"07A5",X"0620",X"05E2",X"05ED",X"0299",X"000E",X"0110",X"00BD",X"FC44",X"F48A",X"F090",X"F1C7",X"F711",X"FED1",X"0754",X"0B1E",X"0932",X"06C5",X"05BC",X"061B",X"04BB",X"010C",X"00C0",X"01A2",X"0022",X"F992",X"F2E9",X"F0BD",X"F335",X"F92C",X"01D7",X"0927",X"0A77",X"0844",X"0666",X"05F5",X"064C",X"0304",X"00BA",X"0137",X"01A9",X"FE12",X"F6D0",X"F1C1",X"F12A",X"F4D8",X"FBFA",X"0501",X"0A33",X"099B",X"076F",X"05C9",X"067D",X"0547",X"01FB",X"011D",X"01D2",X"0128",X"FB81",X"F4AB",X"F0E3",X"F1CC",X"F67D",X"FEFB",X"0793",X"0A6D",X"0947",X"06DC",X"064A",X"06A9",X"0390",X"013F",X"0105",X"0214",X"FF6D",X"F925",X"F35B",X"F166",X"F351",X"F947",X"02AC",X"0921",X"09F8",X"07FA",X"05B7",X"0674",X"0503",X"0215",X"00A3",X"01CA",X"0202",X"FDC4",X"F723",X"F28B",X"F1CF",X"F4A9",X"FC60",X"0587",X"0991",X"0978",X"06C8",X"0647",X"0670",X"03F1",X"0171",X"00F8",X"0293",X"011F",X"FBA1",X"F55E",X"F215",X"F231",X"F68A",X"FFC1",X"072B",X"09D3",X"0854",X"0634",X"06A9",X"0572",X"02E0",X"00E4",X"0202",X"02B3",X"FFA5",X"F952",X"F3F8",X"F1C8",X"F2B3",X"F970",X"02B0",X"0865",X"09C4",X"0735",X"06A7",X"065E",X"0481",X"01BF",X"013D",X"02D1",X"0260",X"FDAF",X"F758",X"F348",X"F18B",X"F426",X"FCB6",X"04B6",X"0966",X"088B",X"06E3",X"06E7",X"05F1",X"0367",X"0119",X"01CA",X"02FF",X"00FC",X"FB61",X"F5EB",X"F2BC",X"F1B4",X"F71F",X"FFD3",X"071C",X"0969",X"0780",X"06D6",X"0681",X"04DA",X"01DB",X"00EB",X"028B",X"030D",X"FF9A",X"F9B9",X"F55A",X"F1F1",X"F2CE",X"F9DE",X"022D",X"0830",X"0833",X"0716",X"06DB",X"0659",X"03CF",X"0162",X"01B3",X"0351",X"025B",X"FD55",X"F82A",X"F3FC",X"F13B",X"F4F8",X"FC94",X"04FD",X"0855",X"0792",X"06F7",X"06FD",X"059F",X"02B5",X"013F",X"0283",X"0393",X"00D4",X"FB6D",X"F71F",X"F26C",X"F1EF",X"F71A",X"FFB2",X"06A8",X"07E6",X"074C",X"0739",X"06FD",X"04AA",X"01F5",X"0199",X"0330",X"0310",X"FEC0",X"FA40",X"F573",X"F1A8",X"F349",X"F9C5",X"02BE",X"0734",X"0794",X"0730",X"0767",X"0654",X"0374",X"0177",X"0216",X"03BA",X"01A8",X"FD08",X"F8C7",X"F373",X"F1A7",X"F4B0",X"FD23",X"04D6",X"0787",X"0779",X"0794",X"078F",X"0598",X"02A3",X"018B",X"030F",X"038C",X"FFB1",X"FBDA",X"F69A",X"F247",X"F1D7",X"F753",X"004A",X"061A",X"0779",X"076E",X"07C2",X"06F6",X"0439",X"01E3",X"01ED",X"03F7",X"024A",X"FEB8",X"FA7B",X"F4F2",X"F1AA",X"F306",X"FA89",X"02B1",X"06C2",X"0758",X"0792",X"07C3",X"060E",X"0313",X"013E",X"02E6",X"03CB",X"00E3",X"FDA7",X"F882",X"F3BB",X"F176",X"F54F",X"FDD4",X"04A7",X"0725",X"0780",X"0800",X"0780",X"04FD",X"01EA",X"017B",X"03AD",X"0253",X"FFBA",X"FBAC",X"F6AB",X"F23D",X"F1E9",X"F83C",X"00C5",X"0606",X"077F",X"0805",X"0848",X"06BA",X"03A3",X"00E0",X"029A",X"0372",X"01BE",X"FEC4",X"FA60",X"F552",X"F193",X"F3B0",X"FB5A",X"02C5",X"0644",X"071E",X"0801",X"07B9",X"05B2",X"020B",X"017D",X"0393",X"0308",X"0110",X"FD7E",X"F8FE",X"F3C6",X"F190",X"F61E",X"FE36",X"0416",X"063B",X"074F",X"07FE",X"0734",X"0423",X"0106",X"0292",X"037F",X"0290",X"0011",X"FC75",X"F76A",X"F28E",X"F28E",X"F8FE",X"009E",X"04E0",X"0677",X"07B3",X"07F3",X"0692",X"0263",X"01AD",X"0347",X"0369",X"01BD",X"FEC5",X"FADA",X"F553",X"F175",X"F424",X"FBAB",X"0254",X"0551",X"072E",X"080B",X"0864",X"0518",X"01DC",X"029A",X"03A5",X"0329",X"00DE",X"FDC6",X"F922",X"F361",X"F193",X"F66C",X"FE37",X"0330",X"05C5",X"0741",X"0859",X"076F",X"033A",X"0208",X"0328",X"03DE",X"026D",X"FFF5",X"FCBE",X"F733",X"F21E",X"F2BA",X"F94C",X"0045",X"0409",X"065C",X"0799",X"08AD",X"058A",X"022B",X"022C",X"0367",X"0376",X"01AE",X"FF55",X"FB54",X"F542",X"F1C8",X"F4CD",X"FC3D",X"01A8",X"0518",X"069A",X"0884",X"07E0",X"03D4",X"01EF",X"0290",X"038A",X"02B8",X"00C9",X"FE68",X"F938",X"F378",X"F1F9",X"F789",X"FE2F",X"0304",X"057D",X"0750",X"08F6",X"0646",X"02F2",X"0229",X"0360",X"03AB",X"0227",X"0058",X"FCE0",X"F6E4",X"F1D0",X"F355",X"F9BE",X"FFB9",X"03FD",X"05E7",X"089D",X"0873",X"04D5",X"023D",X"0272",X"03AE",X"0320",X"017B",X"FFBB",X"FB56",X"F4FF",X"F1EA",X"F5F2",X"FBE8",X"0187",X"0449",X"06E7",X"08F8",X"06EE",X"0351",X"01E5",X"0304",X"03C9",X"0290",X"0144",X"FEB2",X"F947",X"F306",X"F2E6",X"F7B9",X"FDFF",X"026D",X"0501",X"0830",X"0899",X"056C",X"026A",X"0229",X"039B",X"0349",X"021A",X"00B8",X"FD65",X"F6B5",X"F25D",X"F467",X"F9DB",X"FFEB",X"0303",X"063A",X"08F5",X"07AA",X"040B",X"01EF",X"02D3",X"03BA",X"02EC",X"01F0",X"0051",X"FB4A",X"F458",X"F298",X"F5C7",X"FC4E",X"00EF",X"03E7",X"079C",X"08F6",X"066E",X"02FA",X"0212",X"0376",X"0373",X"0288",X"0190",X"FF23",X"F84B",X"F300",X"F2F7",X"F7EB",X"FE0F",X"01A1",X"054F",X"08CC",X"088E",X"0531",X"0253",X"02D8",X"039D",X"031D",X"020C",X"015F",X"FCF0",X"F5F8",X"F28A",X"F468",X"FA90",X"FF62",X"02D8",X"0703",X"0927",X"0762",X"038C",X"0214",X"02FB",X"0345",X"026B",X"020C",X"00A3",X"FA83",X"F4BC",X"F2BC",X"F690",X"FC65",X"002E",X"0423",X"0804",X"08D1",X"05DA",X"027E",X"027B",X"0365",X"033F",X"0244",X"0281",X"FEDB",X"F877",X"F373",X"F3A5",X"F8DB",X"FD94",X"014D",X"05CD",X"08D2",X"081E",X"0413",X"021A",X"029B",X"0362",X"0257",X"028C",X"01B8",X"FCBA",X"F679",X"F2E9",X"F582",X"FAC8",X"FEA0",X"02C9",X"0724",X"091A",X"067C",X"02E8",X"020D",X"032C",X"02F8",X"0246",X"0310",X"0085",X"FACF",X"F4BD",X"F34C",X"F78C",X"FBEC",X"FFC5",X"044A",X"0862",X"089D",X"0509",X"0276",X"0288",X"0373",X"024A",X"02E6",X"02A4",X"FECD",X"F85A",X"F35E",X"F486",X"F909",X"FCE2",X"010C",X"05D9",X"08F8",X"0741",X"03D4",X"0223",X"0354",X"02D5",X"0279",X"036F",X"01F3",X"FD04",X"F648",X"F33D",X"F62B",X"FA31",X"FE01",X"026E",X"076A",X"08AF",X"0610",X"02B6",X"02BA",X"036B",X"027C",X"032C",X"0373",X"00DB",X"FAB3",X"F46F",X"F40B",X"F772",X"FB41",X"FF18",X"0455",X"0870",X"080E",X"048F",X"0261",X"0358",X"02C3",X"026E",X"0355",X"02CC",X"FF05",X"F7E9",X"F3B8",X"F543",X"F8DE",X"FC66",X"00DD",X"0686",X"08F6",X"0710",X"0338",X"02F1",X"0349",X"025E",X"02CA",X"037A",X"0235",X"FCB0",X"F5DD",X"F409",X"F65C",X"F9E8",X"FD6B",X"02FD",X"07BD",X"08AD",X"0523",X"02B5",X"031D",X"028B",X"023D",X"0316",X"0391",X"010E",X"FA10",X"F4E1",X"F4BF",X"F7BB",X"FABD",X"FF2E",X"04E8",X"08AA",X"07A9",X"03D7",X"0322",X"0318",X"0247",X"027A",X"036C",X"035D",X"FEB1",X"F7C1",X"F481",X"F5DA",X"F8BF",X"FBE0",X"0127",X"067A",X"08DA",X"05DE",X"0362",X"035C",X"02B2",X"0241",X"02B6",X"03E2",X"025E",X"FC14",X"F64D",X"F4BE",X"F6F7",X"F961",X"FD73",X"02E8",X"07E0",X"07D4",X"0473",X"036B",X"031B",X"0266",X"024F",X"034A",X"044D",X"0096",X"F9FB",X"F565",X"F5AE",X"F78D",X"FA4D",X"FEEF",X"04FB",X"0887",X"0663",X"03FA",X"038E",X"02E4",X"025D",X"0262",X"040E",X"036C",X"FE1F",X"F7B5",X"F530",X"F652",X"F842",X"FBB6",X"0119",X"071E",X"0836",X"0535",X"03D3",X"0338",X"02A4",X"01E9",X"02CA",X"044F",X"01DC",X"FBBA",X"F673",X"F5C9",X"F6F5",X"F956",X"FD25",X"0380",X"082B",X"06F0",X"0488",X"03A6",X"0318",X"0261",X"01F5",X"03DF",X"0411",X"0007",X"F954",X"F609",X"F60D",X"F786",X"FA09",X"FF04",X"05DE",X"080F",X"05D1",X"043C",X"037C",X"0316",X"01EA",X"02BC",X"046F",X"033E",X"FD7E",X"F7C4",X"F5DA",X"F66F",X"F838",X"FB40",X"01D5",X"076C",X"0740",X"0523",X"03C8",X"0364",X"0253",X"01A1",X"0359",X"048E",X"018D",X"FB09",X"F6FC",X"F5FA",X"F70B",X"F8CE",X"FD3C",X"047A",X"07CD",X"06A1",X"04AF",X"03BF",X"034A",X"01BF",X"0221",X"0418",X"0436",X"FF44",X"F986",X"F691",X"F689",X"F794",X"F9A3",X"FFE1",X"0634",X"0741",X"05A4",X"03DE",X"0381",X"0255",X"0178",X"02CA",X"04D7",X"02EB",X"FD3E",X"F863",X"F689",X"F702",X"F7AD",X"FB58",X"02A5",X"06DF",X"06CD",X"04AB",X"03D9",X"0341",X"01CE",X"01BF",X"03E3",X"04F0",X"0123",X"FB7A",X"F788",X"F6DB",X"F717",X"F818",X"FDFC",X"04A3",X"0723",X"05EE",X"0423",X"03BF",X"0298",X"0162",X"0239",X"04C9",X"03D4",X"FEFE",X"F9B9",X"F71F",X"F722",X"F6E0",X"F9BC",X"00CE",X"0602",X"070F",X"051B",X"042B",X"036D",X"021F",X"015C",X"0374",X"051C",X"0279",X"FD15",X"F872",X"F73C",X"F6CF",X"F6D3",X"FBFD",X"02C7",X"06BA",X"062F",X"04AA",X"0411",X"0335",X"01AE",X"0200",X"049F",X"04AA",X"00B9",X"FB1D",X"F7D3",X"F761",X"F61F",X"F81A",X"FE64",X"049E",X"06B1",X"0564",X"047E",X"03FE",X"02AC",X"014E",X"032B",X"0537",X"03B5",X"FEBA",X"F998",X"F7FA",X"F6C8",X"F603",X"FA0A",X"00E5",X"060A",X"0653",X"0508",X"0465",X"03B4",X"01BC",X"01A1",X"041C",X"0513",X"022D",X"FC79",X"F8BA",X"F7C0",X"F5DF",X"F6E3",X"FC48",X"0339",X"0660",X"05C3",X"04B3",X"0451",X"02F6",X"014A",X"02A5",X"04E5",X"04AF",X"006D",X"FAF5",X"F900",X"F723",X"F5D0",X"F843",X"FED9",X"04A8",X"0619",X"0514",X"0461",X"03E9",X"01F8",X"0169",X"0399",X"054E",X"03BD",X"FE33",X"FA4B",X"F88F",X"F64D",X"F5F7",X"FA41",X"0150",X"0585",X"05D8",X"04B8",X"0481",X"033F",X"0161",X"022E",X"0478",X"0578",X"01DF",X"FC75",X"F9FD",X"F7A1",X"F595",X"F6B8",X"FCCA",X"0337",X"05FB",X"0553",X"04B1",X"0446",X"023F",X"014B",X"0306",X"054D",X"04D4",X"FFA3",X"FBB8",X"F960",X"F6D0",X"F545",X"F869",X"FF30",X"047B",X"05A8",X"04EC",X"04E0",X"03A1",X"0198",X"01CF",X"03EE",X"0605",X"0318",X"FE21",X"FB25",X"F89F",X"F5D3",X"F5A7",X"FAAA",X"0177",X"0544",X"0532",X"04D5",X"0485",X"0286",X"0139",X"0217",X"04FD",X"0567",X"011F",X"FD2A",X"FA8B",X"F7C7",X"F542",X"F716",X"FD52",X"0375",X"057D",X"050F",X"050E",X"03E4",X"01D6",X"012B",X"0328",X"05F7",X"0401",X"FF88",X"FC2C",X"F9A6",X"F665",X"F513",X"F8D4",X"FFB3",X"0481",X"0532",X"050E",X"04DE",X"02F9",X"0161",X"016E",X"04AA",X"05C6",X"026A",X"FE6B",X"FBB8",X"F8C4",X"F594",X"F5F4",X"FB4A",X"01E7",X"04FB",X"0502",X"0537",X"0413",X"022C",X"00B7",X"0267",X"05A7",X"04CE",X"00F7",X"FD90",X"FB1A",X"F77E",X"F512",X"F758",X"FDD9",X"0370",X"04CF",X"0532",X"04F8",X"036D",X"0144",X"0094",X"03C8",X"05A5",X"036C",X"FFAD",X"FD11",X"FA0B",X"F66C",X"F565",X"F98A",X"0050",X"0421",X"04E4",X"0547",X"0469",X"02BD",X"0081",X"01B1",X"0512",X"054D",X"0214",X"FEC3",X"FC3B",X"F89B",X"F54E",X"F605",X"FBD9",X"020C",X"0435",X"053A",X"0518",X"0436",X"01D2",X"007E",X"0320",X"05B3",X"045E",X"00D2",X"FE20",X"FB32",X"F732",X"F4D2",X"F784",X"FE5E",X"02D0",X"04A1",X"053E",X"0509",X"0395",X"00CC",X"0147",X"047E",X"0594",X"02EE",X"FFD8",X"FD69",X"F9F7",X"F5FC",X"F511",X"FA18",X"0049",X"038C",X"0508",X"053B",X"04E3",X"0242",X"0052",X"023C",X"0548",X"04B5",X"01B3",X"FF22",X"FC8D",X"F893",X"F4F7",X"F654",X"FC94",X"018E",X"0438",X"0504",X"0551",X"041B",X"0120",X"00A5",X"03AF",X"0595",X"03BD",X"00D3",X"FE96",X"FB72",X"F70C",X"F47F",X"F871",X"FE69",X"028D",X"046A",X"051A",X"0544",X"02EB",X"0075",X"01A2",X"04DC",X"053D",X"02A1",X"004D",X"FDEE",X"FA43",X"F57B",X"F560",X"FAA0",X"FFF7",X"034E",X"0467",X"0560",X"04AE",X"0191",X"0031",X"02D5",X"054B",X"0434",X"01C8",X"FFBA",X"FD20",X"F88E",X"F4DE",X"F74D",X"FCA8",X"0174",X"03A7",X"04C4",X"056C",X"0382",X"0081",X"00E8",X"0424",X"0529",X"0346",X"0126",X"FF1F",X"FBDE",X"F685",X"F52F",X"F8F4",X"FE7E",X"0249",X"03D6",X"0539",X"0519",X"022B",X"0044",X"023F",X"050C",X"0490",X"027D",X"0069",X"FE68",X"F9BF",X"F54F",X"F61A",X"FAD1",X"0019",X"02DF",X"0490",X"05C6",X"044A",X"010E",X"009A",X"03A4",X"0528",X"03E5",X"01B2",X"0015",X"FD3F",X"F7B3",X"F521",X"F76B",X"FCCB",X"0108",X"032B",X"050B",X"0584",X"02E8",X"0051",X"01A8",X"0484",X"04DC",X"0325",X"0137",X"FFCC",X"FB3E",X"F654",X"F587",X"F952",X"FE98",X"01C7",X"03C3",X"0576",X"04B6",X"01A0",X"0077",X"02F7",X"04E4",X"0467",X"023A",X"0123",X"FE96",X"F93C",X"F586",X"F670",X"FB45",X"FFEB",X"0252",X"048D",X"05A5",X"03AF",X"00B9",X"0158",X"03E4",X"04F6",X"0379",X"01BA",X"00BB",X"FCAF",X"F786",X"F53F",X"F7E6",X"FD3B",X"00B9",X"031B",X"053B",X"0550",X"022F",X"0076",X"0241",X"048B",X"04A7",X"0289",X"01DE",X"FFC8",X"FAF3",X"F652",X"F5C3",X"F9DF",X"FE89",X"0151",X"03D2",X"05B3",X"043A",X"0102",X"00DE",X"0331",X"050B",X"03B8",X"025F",X"01B3",X"FE82",X"F93D",X"F59C",X"F6FF",X"FBCA",X"FF85",X"0211",X"04B5",X"0588",X"0297",X"007C",X"0176",X"041D",X"0497",X"02E6",X"0263",X"00F0",X"FCCF",X"F7B3",X"F5A9",X"F8CF",X"FD36",X"0051",X"02FE",X"0587",X"0491",X"0183",X"0097",X"0297",X"04D3",X"03ED",X"02CF",X"024C",X"FFD8",X"FAE0",X"F63A",X"F64E",X"FA49",X"FE44",X"00FA",X"040B",X"059F",X"0347",X"00EB",X"0119",X"03DB",X"04AC",X"0372",X"02F7",X"01FE",X"FE73",X"F8FD",X"F5A1",X"F782",X"FBBB",X"FF0A",X"01E6",X"050A",X"04C7",X"022A",X"0069",X"0205",X"047D",X"042E",X"0337",X"02F7",X"0133",X"FCB8",X"F745",X"F5F3",X"F919",X"FD24",X"FFDD",X"035F",X"0565",X"03E4",X"0131",X"0091",X"031E",X"046B",X"0393",X"0325",X"029B",X"0000",X"FA7E",X"F64C",X"F6EF",X"FAE9",X"FE06",X"0109",X"048F",X"0510",X"02CF",X"005E",X"016D",X"03EC",X"0404",X"0360",X"0318",X"0224",X"FE31",X"F88B",X"F5F6",X"F839",X"FC09",X"FECA",X"0297",X"052E",X"04A5",X"01A8",X"006A",X"028A",X"0417",X"03AC",X"032F",X"0305",X"014B",X"FC1E",X"F717",X"F661",X"F9C3",X"FCB4",X"000A",X"03D0",X"0560",X"0390",X"009D",X"0106",X"0351",X"03E2",X"0368",X"033A",X"0303",X"FFD6",X"FA2D",X"F655",X"F7AA",X"FAE7",X"FDA5",X"0176",X"04A7",X"0503",X"0225",X"0045",X"01F6",X"03AB",X"03B8",X"033E",X"037E",X"028E",X"FE25",X"F865",X"F66C",X"F8E3",X"FB89",X"FECB",X"02A0",X"0507",X"03EA",X"00D9",X"00AC",X"02C5",X"03D9",X"039E",X"0384",X"03D5",X"0183",X"FC15",X"F708",X"F735",X"F9B2",X"FC7D",X"0018",X"03CA",X"0513",X"02A2",X"0056",X"016B",X"032D",X"03B4",X"0346",X"03C9",X"037F",X"0011",X"F9EE",X"F6D4",X"F818",X"FA76",X"FD99",X"016E",X"04A2",X"045A",X"0145",X"0083",X"021E",X"03A5",X"0371",X"0388",X"0417",X"02F8",X"FDEE",X"F844",X"F724",X"F8B7",X"FB49",X"FEB2",X"02AC",X"04FD",X"031D",X"00B4",X"010F",X"02DC",X"03AA",X"0361",X"03D2",X"0435",X"01AC",X"FB78",X"F789",X"F78C",X"F97B",X"FC2D",X"FFF2",X"03F1",X"0497",X"01F4",X"009D",X"01C7",X"0363",X"036E",X"0372",X"040B",X"03FC",X"FF8F",X"F9BF",X"F769",X"F839",X"FA67",X"FD6C",X"01AE",X"04D3",X"03AA",X"0135",X"00B7",X"025D",X"033F",X"032B",X"036B",X"0478",X"02F1",X"FD40",X"F899",X"F7A7",X"F8DB",X"FB32",X"FEAC",X"0346",X"04BC",X"02A5",X"00B6",X"0149",X"02D3",X"0334",X"030E",X"03BE",X"0492",X"011C",X"FB59",X"F81A",X"F7FB",X"F9AB",X"FC2D",X"0091",X"044C",X"0418",X"01B5",X"009D",X"01E8",X"02E3",X"0300",X"02FF",X"048B",X"0410",X"FF26",X"FA28",X"F7F2",X"F87E",X"FA33",X"FD4F",X"0228",X"045D",X"030E",X"00D4",X"00F6",X"0239",X"0309",X"02B7",X"038F",X"050E",X"02A7",X"FD45",X"F930",X"F81A",X"F911",X"FADF",X"FF22",X"035C",X"043C",X"0209",X"00B0",X"016D",X"02BA",X"0301",X"02CD",X"0490",X"04E4",X"00CD",X"FB8E",X"F861",X"F844",X"F921",X"FBCE",X"00BA",X"0402",X"0387",X"0159",X"00EB",X"01FF",X"02FF",X"028D",X"0347",X"053E",X"03BF",X"FEF6",X"FA3D",X"F866",X"F89D",X"F9B6",X"FD9E",X"0247",X"0430",X"027C",X"0100",X"0130",X"0293",X"02EA",X"028F",X"043F",X"0550",X"0277",X"FD45",X"F963",X"F88C",X"F89B",X"FAB9",X"FF3B",X"0348",X"0384",X"01A1",X"00A6",X"019B",X"02D1",X"0250",X"02CA",X"0509",X"04B1",X"00B8",X"FBA7",X"F920",X"F885",X"F917",X"FC42",X"0112",X"03C3",X"02EB",X"0131",X"00DE",X"024F",X"02AF",X"0221",X"03C3",X"055C",X"03A4",X"FED6",X"FA93",X"F8FB",X"F87A",X"F9D9",X"FDF6",X"0279",X"038D",X"021B",X"00A8",X"013F",X"029C",X"022B",X"027E",X"049E",X"052A",X"022E",X"FCFB",X"FA02",X"F8A1",X"F892",X"FAF1",X"FFE6",X"032D",X"032E",X"0169",X"0094",X"01FD",X"0287",X"01E9",X"0347",X"0526",X"04B8",X"004C",X"FBF3",X"F99D",X"F886",X"F8FC",X"FCA8",X"0159",X"0380",X"0289",X"00B0",X"00EB",X"027B",X"0206",X"0221",X"03FD",X"0589",X"0356",X"FEAB",X"FB27",X"F930",X"F857",X"F9DF",X"FE65",X"0246",X"0341",X"01A8",X"005C",X"01B3",X"0269",X"01E8",X"02D5",X"04FE",X"057A",X"01CB",X"FD77",X"FA86",X"F8D1",X"F867",X"FB59",X"FFE9",X"02D3",X"02AD",X"00C4",X"00BD",X"0246",X"0217",X"0207",X"037B",X"05BB",X"0456",X"000B",X"FC38",X"F9F4",X"F84D",X"F902",X"FCF3",X"0126",X"0306",X"01D9",X"0069",X"0199",X"025E",X"01DC",X"0229",X"0484",X"0594",X"02D3",X"FE94",X"FB7F",X"F961",X"F855",X"FA75",X"FECB",X"024E",X"02F4",X"00E6",X"00AD",X"01E3",X"0200",X"019E",X"02DF",X"056B",X"04FF",X"016F",X"FD81",X"FAD4",X"F8AD",X"F8AD",X"FBD0",X"000A",X"02E2",X"0218",X"0073",X"013C",X"0215",X"01DD",X"01B5",X"03F2",X"05AE",X"03F0",X"FFF8",X"FCAC",X"FA0D",X"F85C",X"F992",X"FD42",X"0167",X"02EC",X"012E",X"00A0",X"0187",X"0208",X"0153",X"0249",X"04E0",X"0575",X"028E",X"FED9",X"FBE1",X"F940",X"F86B",X"FA95",X"FEB8",X"0277",X"024B",X"00CC",X"00FC",X"020C",X"01D8",X"0170",X"0356",X"0594",X"04B4",X"0130",X"FDD8",X"FAD8",X"F883",X"F8BD",X"FBB0",X"0053",X"02AD",X"0187",X"00B3",X"0174",X"022C",X"016B",X"01EA",X"0471",X"05B9",X"03A4",X"0014",X"FCDF",X"F9C5",X"F84A",X"F974",X"FD42",X"0198",X"0245",X"0102",X"00C3",X"01E2",X"01D3",X"013D",X"02AE",X"0550",X"0562",X"0286",X"FF42",X"FBF8",X"F91B",X"F874",X"FA6B",X"FF28",X"021E",X"01B2",X"008D",X"0114",X"01EE",X"014D",X"015E",X"03BA",X"05B3",X"0469",X"016A",X"FE25",X"FAB5",X"F8B4",X"F8B7",X"FC17",X"00AF",X"0252",X"0148",X"00B2",X"01AE",X"01CD",X"010A",X"0202",X"04D9",X"0588",X"0367",X"0078",X"FCEC",X"F9E9",X"F85A",X"F969",X"FDE2",X"0182",X"01DD",X"00AC",X"00F3",X"01E2",X"0170",X"0101",X"0316",X"057B",X"0503",X"028E",X"FF52",X"FBB2",X"F93A",X"F827",X"FACD",X"FF69",X"01E7",X"0148",X"0095",X"0179",X"01E5",X"00FA",X"0199",X"0451",X"05B1",X"043C",X"01B1",X"FE04",X"FAE3",X"F888",X"F8CB",X"FC91",X"00C9",X"01EC",X"00C9",X"00C4",X"01B3",X"0158",X"00A0",X"0240",X"04DF",X"050F",X"036C",X"0068",X"FCF7",X"FA11",X"F84B",X"FA0D",X"FE7E",X"01BF",X"018E",X"00A0",X"0136",X"01B4",X"00C4",X"00DA",X"0365",X"0521",X"04AE",X"029F",X"FF43",X"FC16",X"F91D",X"F873",X"FB61",X"FFE5",X"01D4",X"0110",X"00BC",X"01A6",X"016D",X"0078",X"01A7",X"043D",X"0520",X"0463",X"0198",X"FE4C",X"FAF9",X"F873",X"F900",X"FCF7",X"00D3",X"0173",X"0089",X"00F9",X"01B9",X"00E9",X"0080",X"02BE",X"04B6",X"054B",X"03A3",X"00A1",X"FD73",X"FA08",X"F847",X"FA3A",X"FE9E",X"0142",X"00F2",X"0089",X"0151",X"0172",X"0056",X"013C",X"0380",X"0501",X"04E5",X"029B",X"FFA6",X"FC4F",X"F93E",X"F89B",X"FBBD",X"FFD6",X"013C",X"0081",X"00C2",X"01B0",X"00F4",X"004E",X"021E",X"041C",X"054C",X"0439",X"01A3",X"FE8C",X"FB0B",X"F871",X"F945",X"FD56",X"00B5",X"00FD",X"008C",X"0163",X"01B4",X"0069",X"00FA",X"02D1",X"04B7",X"0522",X"0360",X"00BC",X"FD6D",X"F9DC",X"F83E",X"FA7A",X"FEB2",X"00C8",X"007C",X"0097",X"01B3",X"0106",X"006B",X"0198",X"0394",X"053F",X"04CF",X"02C5",X"FFE7",X"FC5A",X"F906",X"F8AB",X"FC13",X"FFD0",X"00B7",X"002E",X"010E",X"0177",X"005E",X"0084",X"0200",X"0437",X"0536",X"0443",X"01E7",X"FEE5",X"FB22",X"F893",X"F9AF",X"FDC1",X"0085",X"007C",X"0081",X"0196",X"00F8",X"0038",X"00BE",X"02A4",X"04A8",X"0508",X"0382",X"0107",X"FDAC",X"F9E1",X"F86B",X"FB24",X"FF10",X"009E",X"0029",X"0111",X"0165",X"0096",X"0050",X"0158",X"0393",X"051B",X"04BC",X"02DD",X"001B",X"FC51",X"F8D5",X"F8F8",X"FC6D",X"FFBF",X"001A",X"0058",X"015E",X"0110",X"0068",X"0088",X"0225",X"0458",X"053E",X"0440",X"0219",X"FF01",X"FAFB",X"F894",X"FA1D",X"FE0F",X"0016",X"FFFD",X"00C9",X"012B",X"0091",X"0000",X"00C0",X"02CF",X"04BE",X"04FE",X"03AD",X"015E",X"FDD2",X"F9DB",X"F8BF",X"FB93",X"FF18",X"FFD8",X"0042",X"0116",X"0113",X"0069",X"0034",X"016A",X"03AE",X"04FC",X"049A",X"02DA",X"0042",X"FC2B",X"F8F7",X"F94D",X"FD20",X"FF72",X"FFCE",X"00B3",X"0147",X"0100",X"005A",X"008B",X"0242",X"0456",X"0516",X"0414",X"023B",X"FEFD",X"FACB",X"F881",X"FA94",X"FE3A",X"FF5C",X"0007",X"00DD",X"0115",X"0098",X"0034",X"00F6",X"0301",X"04B7",X"04C3",X"038F",X"0152",X"FD8F",X"F9B1",X"F8F1",X"FC42",X"FED0",X"FF93",X"0062",X"0117",X"0100",X"0064",X"0038",X"0199",X"03AD",X"04EB",X"046A",X"0303",X"0045",X"FC2F",X"F8DC",X"FA22",X"FD69",X"FF13",X"FFE2",X"00AE",X"00E6",X"00AF",X"0010",X"0068",X"0233",X"044A",X"04C4",X"0415",X"0241",X"FF04",X"FAA1",X"F8E0",X"FB6C",X"FE12",X"FF51",X"0035",X"00CB",X"00EE",X"0074",X"002D",X"010A",X"0333",X"04BB",X"04CC",X"03BC",X"017F",X"FD84",X"F963",X"F992",X"FC52",X"FE59",X"FF78",X"004E",X"00B6",X"00B0",X"0017",X"0029",X"01B1",X"03E8",X"04EE",X"04A3",X"0337",X"008C",X"FBBE",X"F90F",X"FA93",X"FD28",X"FEB8",X"FFC5",X"0069",X"00CB",X"007A",X"0009",X"007E",X"029F",X"0464",X"04F4",X"0446",X"02BE",X"FF03",X"FA50",X"F967",X"FBA1",X"FDC7",X"FF2F",X"000B",X"00A8",X"00A5",X"0037",X"FFE7",X"0113",X"0339",X"04BD",X"04BF",X"03DD",X"01CB",X"FD08",X"F96D",X"F9FD",X"FC52",X"FE34",X"FF66",X"0038",X"00B5",X"00B5",X"0030",X"0046",X"01EF",X"03E6",X"04DD",X"046F",X"0399",X"0049",X"FB5D",X"F970",X"FAED",X"FD0B",X"FEB5",X"FFCD",X"0086",X"00C8",X"0071",X"FFDF",X"009E",X"027E",X"0459",X"04A3",X"0462",X"02E8",X"FE7D",X"FA4B",X"F9DE",X"FB9C",X"FDA3",X"FF11",X"001A",X"0086",X"00A6",X"0002",X"FFE5",X"011C",X"0354",X"048B",X"0493",X"0461",X"01C2",X"FCB8",X"F9FC",X"FA81",X"FC79",X"FE2E",X"FF87",X"003E",X"00A6",X"006C",X"FFC0",X"0014",X"01D1",X"03E6",X"0465",X"049E",X"03E5",X"FFEB",X"FB60",X"F9E7",X"FB28",X"FD1A",X"FEC6",X"FFE6",X"0082",X"00C1",X"001A",X"FFBC",X"0075",X"02B0",X"041B",X"0460",X"04D5",X"02E4",X"FE30",X"FAB4",X"FA55",X"FBEE",X"FDBB",X"FF47",X"0000",X"008B",X"005A",X"FFC4",X"FF9B",X"012E",X"0367",X"0432",X"04B5",X"04A7",X"0142",X"FCAA",X"FA41",X"FAD5",X"FC89",X"FE5E",X"FF8A",X"0049",X"008F",X"0026",X"FF78",X"FFDE",X"0219",X"03AC",X"0441",X"0525",X"03F7",X"FFA8",X"FBA9",X"FA71",X"FB5B",X"FD3B",X"FED2",X"FFC5",X"0063",X"005F",X"FFE5",X"FF55",X"0099",X"02D7",X"03CF",X"04C5",X"052E",X"0294",X"FDF7",X"FACD",X"FA7E",X"FBD8",X"FDC9",X"FF19",X"0013",X"0072",X"005D",X"FF87",X"FF89",X"0190",X"0345",X"0401",X"0543",X"04B4",X"010C",X"FCAA",X"FA94",X"FADA",X"FC99",X"FE49",X"FF88",X"002D",X"0083",X"0014",X"FF39",X"0015",X"024F",X"0350",X"0476",X"055F",X"03A8",X"FF57",X"FBBC",X"FA7F",X"FB5E",X"FD30",X"FEB3",X"FFC5",X"0053",X"0088",X"FFA5",X"FF45",X"0112",X"02B8",X"0396",X"0505",X"0538",X"0241",X"FDEA",X"FB11",X"FA97",X"FC05",X"FDBF",X"FF34",X"FFF3",X"007C",X"0045",X"FF39",X"FFBE",X"01BB",X"02DA",X"0414",X"056A",X"047B",X"00B3",X"FCD2",X"FAA3",X"FB0D",X"FC9F",X"FE5F",X"FF7F",X"0022",X"009C",X"FFD3",X"FF0B",X"007B",X"0204",X"031D",X"04AC",X"0598",X"0370",X"FF6E",X"FBF6",X"FABD",X"FB80",X"FD31",X"FED7",X"FFB1",X"006B",X"007D",X"FF39",X"FF6D",X"010A",X"022E",X"0356",X"051E",X"050F",X"0212",X"FE19",X"FB54",X"FAE5",X"FC07",X"FDDE",X"FF25",X"FFE8",X"00C1",X"FFFF",X"FF06",X"0011",X"0194",X"028A",X"0423",X"059B",X"0448",X"00C9",X"FCF9",X"FB06",X"FB20",X"FC8E",X"FE3F",X"FF2C",X"003E",X"00A7",X"FF5F",X"FF5F",X"00C0",X"01D7",X"0311",X"04FB",X"0564",X"033A",X"FF4F",X"FC21",X"FADD",X"FB89",X"FD42",X"FE90",X"FF86",X"00A2",X"001A",X"FF20",X"FFBA",X"010F",X"01F3",X"03AD",X"055D",X"04F0",X"0209",X"FE32",X"FB9F",X"FB0E",X"FC42",X"FDF0",X"FED6",X"001F",X"009D",X"FF77",X"FF22",X"003E",X"013C",X"025A",X"0471",X"0578",X"042A",X"00B4",X"FD22",X"FB2D",X"FB50",X"FCF5",X"FE28",X"FF2F",X"0094",X"001C",X"FF11",X"FF7C",X"00B2",X"016A",X"031E",X"0502",X"0562",X"0318",X"FF64",X"FC46",X"FAF7",X"FBD8",X"FD79",X"FE54",X"FFCB",X"009B",X"FFAC",X"FF04",X"0000",X"00D5",X"01E7",X"03D6",X"0560",X"04D0",X"01E6",X"FE4D",X"FBAD",X"FB29",X"FC9D",X"FDAA",X"FECA",X"004A",X"0038",X"FEFB",X"FF3E",X"0032",X"010C",X"0288",X"0494",X"0589",X"0413",X"00BB",X"FD53",X"FB38",X"FBB2",X"FD0E",X"FDE9",X"FF6F",X"007F",X"FFAB",X"FEFC",X"FFB5",X"006F",X"016D",X"0339",X"0517",X"054B",X"0309",X"FF93",X"FC66",X"FB34",X"FC48",X"FD2C",X"FE4C",X"FFEA",X"0045",X"FF1C",X"FF2B",X"FFF1",X"00B6",X"01F4",X"03F5",X"0571",X"04B6",X"01F7",X"FE7F",X"FBA8",X"FBA4",X"FCA7",X"FD7B",X"FEE8",X"0058",X"FFC2",X"FF00",X"FF68",X"0027",X"00F2",X"029C",X"04AB",X"057A",X"03E7",X"00F7",X"FD42",X"FB8D",X"FC22",X"FCEE",X"FDDD",X"FF95",X"0026",X"FF34",X"FEF8",X"FF90",X"003E",X"0156",X"0355",X"052C",X"050F",X"0327",X"FFAB",X"FC57",X"FBB4",X"FC6C",X"FD20",X"FE88",X"0019",X"FFBF",X"FEF4",X"FF27",X"FFDF",X"0090",X"0208",X"0437",X"0575",X"04A4",X"0227",X"FE4B",X"FBE5",X"FBF1",X"FC9C",X"FD61",X"FF54",X"001C",X"FF58",X"FEF0",X"FF69",X"FFF8",X"00D0",X"02AE",X"04D5",X"053A",X"0417",X"00D3",X"FD2D",X"FBBD",X"FC38",X"FC99",X"FE02",X"FFC4",X"FFD9",X"FF17",X"FF1B",X"FFA2",X"0032",X"015D",X"039E",X"052C",X"052D",X"0353",X"FF70",X"FC78",X"FC01",X"FC3B",X"FCCB",X"FEC6",X"0003",X"FF90",X"FF00",X"FF3E",X"FFC2",X"0053",X"0206",X"043A",X"052B",X"04D7",X"020B",X"FE28",X"FC30",X"FC2F",X"FC31",X"FD8D",X"FF70",X"FFEB",X"FF3A",X"FF05",X"FF66",X"FFE1",X"00CB",X"02F5",X"0497",X"0555",X"042F",X"00AC",X"FD3C",X"FC49",X"FC17",X"FC84",X"FE5D",X"FFD1",X"FF97",X"FF07",X"FF1D",X"FF9C",X"FFED",X"017E",X"038E",X"04F7",X"053D",X"0321",X"FF30",X"FCCB",X"FC2D",X"FC00",X"FD1E",X"FF1B",X"FFD6",X"FF61",X"FEFB",X"FF65",X"FF89",X"004A",X"0241",X"0402",X"053E",X"04E8",X"01C5",X"FE2D",X"FCB5",X"FC18",X"FC4A",X"FDF6",X"FF8B",X"FFA7",X"FEFE",X"FEFA",X"FF4B",X"FF82",X"00F7",X"02DC",X"0476",X"0565",X"041A",X"0054",X"FD99",X"FC8C",X"FC1E",X"FCE3",X"FEC1",X"FFBE",X"FF6F",X"FEC5",X"FF14",X"FF1A",X"FFDC",X"019D",X"0360",X"04D8",X"0571",X"02D9",X"FF27",X"FD46",X"FC5E",X"FC2A",X"FD87",X"FF3C",X"FFCB",X"FF16",X"FEFB",X"FF18",X"FF39",X"0073",X"023C",X"03ED",X"0571",X"04D0",X"0150",X"FE50",X"FCD9",X"FBFF",X"FC78",X"FE2E",X"FF98",X"FF7C",X"FEFE",X"FF0F",X"FEF8",X"FF96",X"0123",X"02C3",X"0490",X"05C1",X"03C9",X"003F",X"FDE5",X"FC7E",X"FBF0",X"FD00",X"FEC0",X"FFA0",X"FF1E",X"FF10",X"FEFE",X"FEF7",X"0014",X"01A8",X"033F",X"054C",X"056F",X"0286",X"FF51",X"FD74",X"FC24",X"FC3D",X"FDA5",X"FF5C",X"FF6B",X"FF0B",X"FF04",X"FEDA",X"FF3E",X"00A4",X"01FD",X"03F5",X"05AF",X"049A",X"0141",X"FEB2",X"FCDD",X"FBFE",X"FC90",X"FE73",X"FF7E",X"FF56",X"FF30",X"FEFE",X"FEDD",X"FFBB",X"0116",X"0283",X"04CF",X"05A9",X"0361",X"0052",X"FE01",X"FC6A",X"FC00",X"FD35",X"FF08",X"FF5D",X"FF36",X"FF10",X"FEC9",X"FF07",X"0038",X"014D",X"0357",X"0577",X"0526",X"0264",X"FFA1",X"FD70",X"FC28",X"FC2E",X"FDFF",X"FF4E",X"FF5F",X"FF37",X"FEF7",X"FE92",X"FF5F",X"0071",X"01B8",X"0427",X"05CB",X"043E",X"017A",X"FED4",X"FCEE",X"FBE8",X"FCD8",X"FEA5",X"FF59",X"FF53",X"FF2F",X"FE97",X"FEBB",X"FFDA",X"00C3",X"0280",X"051D",X"056B",X"035C",X"008C",X"FE2A",X"FC78",X"FC18",X"FD91",X"FF07",X"FF46",X"FF4D",X"FEF1",X"FE6E",X"FF17",X"000A",X"011D",X"037F",X"0585",X"04E9",X"0274",X"FFB9",X"FD7D",X"FBF4",X"FC6E",X"FE35",X"FF24",X"FF4C",X"FF51",X"FE9A",X"FE9C",X"FF7E",X"002F",X"01BB",X"048B",X"0591",X"043B",X"018E",X"FF19",X"FCDF",X"FBFE",X"FD2D",X"FEB2",X"FF23",X"FF76",X"FEFC",X"FE5C",X"FEE2",X"FFC8",X"0072",X"02D1",X"052D",X"0558",X"0349",X"00B1",X"FE48",X"FC3D",X"FC31",X"FDC2",X"FEB7",X"FF3B",X"FF5D",X"FE9E",X"FE71",X"FF64",X"FFC5",X"012B",X"03C4",X"0577",X"04D4",X"027A",X"FFFD",X"FD6F",X"FC06",X"FCD1",X"FE42",X"FEE7",X"FF74",X"FF0B",X"FE44",X"FEC8",X"FF6F",X"FFEC",X"0203",X"0477",X"0576",X"0407",X"01CC",X"FF2B",X"FCC0",X"FC38",X"FD85",X"FE7C",X"FF44",X"FF81",X"FE9F",X"FE4F",X"FF1A",X"FF59",X"0066",X"02C0",X"0514",X"050D",X"0353",X"0105",X"FE3C",X"FC5A",X"FCBF",X"FDF0",X"FED3",X"FF8F",X"FF40",X"FE3F",X"FEAB",X"FF2B",X"FF7E",X"0108",X"03B1",X"053A",X"0476",X"0298",X"001C",X"FD52",X"FC4D",X"FD34",X"FE32",X"FF1B",X"FFB3",X"FECB",X"FE4D",X"FEFA",X"FF26",X"FFD0",X"01EF",X"048A",X"0518",X"03EF",X"01EE",X"FF1B",X"FCB6",X"FC97",X"FD81",X"FE79",X"FF80",X"FF62",X"FE57",X"FEA6",X"FF12",X"FF3D",X"0052",X"02FD",X"04F0",X"04BC",X"034E",X"010A",X"FDFF",X"FC81",X"FCFC",X"FDDD",X"FEF1",X"FFCA",X"FEDF",X"FE68",X"FED5",X"FF10",X"FF4B",X"012A",X"03CD",X"04F3",X"044C",X"02BA",X"FFE0",X"FD3B",X"FCA7",X"FD4F",X"FE1E",X"FF88",X"FF90",X"FE92",X"FE93",X"FF15",X"FF14",X"FFC7",X"021F",X"045A",X"04BF",X"03E0",X"01E1",X"FEC5",X"FCF5",X"FD05",X"FD7C",X"FEA9",X"FFC0",X"FEFE",X"FE7A",X"FEBC",X"FF08",X"FF08",X"0068",X"0305",X"04A1",X"048A",X"0386",X"00D8",X"FDF3",X"FCEC",X"FD1D",X"FDBD",X"FF49",X"FF77",X"FEAB",X"FE6E",X"FEF3",X"FEE0",X"FF41",X"014D",X"03C6",X"0498",X"0463",X"02C4",X"FFC3",X"FD87",X"FD27",X"FD30",X"FE7F",X"FFA4",X"FF32",X"FE54",X"FE96",X"FEE0",X"FEC1",X"FFC0",X"0242",X"0415",X"049A",X"041D",X"01CF",X"FEB7",X"FD71",X"FD17",X"FD90",X"FF1E",X"FF93",X"FED8",X"FE61",X"FECF",X"FECC",X"FEDB",X"0093",X"0309",X"044B",X"049F",X"0387",X"0090",X"FE19",X"FD47",X"FCF8",X"FE15",X"FF59",X"FF51",X"FE6F",X"FE8F",X"FEE6",X"FEC3",X"FF4F",X"0196",X"0385",X"048A",X"0495",X"02B0",X"FF8B",X"FDF0",X"FD0D",X"FD35",X"FEA0",X"FF81",X"FED3",X"FE4B",X"FEAA",X"FED0",X"FE9B",X"0019",X"025B",X"03EF",X"04BF",X"044C",X"0191",X"FF0F",X"FDAE",X"FCF3",X"FDC4",X"FF2F",X"FF46",X"FE5E",X"FE4F",X"FEAD",X"FE77",X"FEDB",X"00D4",X"02E6",X"042D",X"04E9",X"037D",X"0089",X"FE9E",X"FD3A",X"FD1E",X"FE6B",X"FF7E",X"FF01",X"FE61",X"FE97",X"FEBC",X"FE64",X"FF86",X"01A5",X"034C",X"0496",X"04BC",X"0248",X"FFCE",X"FDF6",X"FCFF",X"FD74",X"FEFC",X"FF68",X"FE98",X"FE3B",X"FEAE",X"FE5D",X"FE93",X"0059",X"025A",X"03C5",X"0522",X"040A",X"0161",X"FF30",X"FD92",X"FCEC",X"FE07",X"FF4B",X"FF19",X"FE4E",X"FE7C",X"FE9D",X"FE3B",X"FF06",X"010A",X"0299",X"0460",X"04FC",X"0318",X"00AB",X"FEAD",X"FD44",X"FD63",X"FECC",X"FF7E",X"FECF",X"FE46",X"FE92",X"FE49",X"FE2E",X"FF98",X"0169",X"0306",X"04EB",X"0465",X"0244",X"0007",X"FE26",X"FD21",X"FDED",X"FF4D",X"FF66",X"FE8B",X"FE88",X"FE8C",X"FE0C",X"FE83",X"0044",X"01C2",X"03EF",X"04F8",X"03AD",X"0179",X"FF59",X"FD87",X"FD39",X"FE6D",X"FF89",X"FEFA",X"FE87",X"FEA5",X"FE67",X"FE17",X"FF5A",X"00BD",X"0283",X"048D",X"04BC",X"02FF",X"00C7",X"FE9E",X"FD23",X"FD79",X"FF01",X"FF4B",X"FE94",X"FE61",X"FE80",X"FDFB",X"FE6F",X"FFCC",X"011C",X"0370",X"04FB",X"0461",X"0250",X"0033",X"FE17",X"FD27",X"FE23",X"FF64",X"FF0E",X"FE75",X"FE8F",X"FE42",X"FDD1",X"FEF0",X"0004",X"01D5",X"0419",X"04E1",X"03A2",X"019F",X"FF58",X"FD86",X"FD57",X"FED4",X"FF6B",X"FECC",X"FE96",X"FEB0",X"FDE2",X"FE4B",X"FF41",X"0069",X"0299",X"0498",X"0482",X"0305",X"00D5",X"FE90",X"FD18",X"FDDF",X"FF39",X"FF3E",X"FEA7",X"FECF",X"FE55",X"FDF7",X"FEBB",X"FF88",X"0112",X"0382",X"04C7",X"0418",X"0258",X"0025",X"FDDD",X"FD2E",X"FE64",X"FF4D",X"FEDB",X"FEAC",X"FEB1",X"FDE3",X"FE2D",X"FEE8",X"FFD1",X"01DF",X"042E",X"04BB",X"03AA",X"01C3",X"FF64",X"FD72",X"FDBA",X"FF06",X"FF3E",X"FEAC",X"FEE6",X"FE44",X"FDDF",X"FE6C",X"FF0A",X"004B",X"02C8",X"0482",X"0471",X"030A",X"0108",X"FE64",X"FD49",X"FE34",X"FF4C",X"FEDA",X"FEEF",X"FEB8",X"FDF9",X"FE1C",X"FEAA",X"FF40",X"0124",X"0370",X"0496",X"03FD",X"0283",X"0015",X"FDC0",X"FD81",X"FECB",X"FF23",X"FEE1",X"FF12",X"FE73",X"FE01",X"FE5F",X"FEC1",X"FFB9",X"01F8",X"040B",X"0483",X"039A",X"01CD",X"FF23",X"FD73",X"FDF6",X"FF17",X"FEE9",X"FF03",X"FED6",X"FE14",X"FE08",X"FE6B",X"FEC6",X"005F",X"02C1",X"0462",X"0454",X"034D",X"0102",X"FE62",X"FD72",X"FEA6",X"FF05",X"FEF3",X"FF0D",X"FE72",X"FDEE",X"FE42",X"FE69",X"FF2F",X"012A",X"037D",X"045E",X"042A",X"02A8",X"0000",X"FDBB",X"FDF5",X"FEF6",X"FEE9",X"FF24",X"FEED",X"FE22",X"FE17",X"FE57",X"FE7D",X"FFA1",X"0208",X"03E5",X"0464",X"03CE",X"01D5",X"FEE9",X"FD8A",X"FE77",X"FEE1",X"FF13",X"FF45",X"FE99",X"FE00",X"FE30",X"FE43",X"FEB2",X"006B",X"02DD",X"0428",X"0479",X"0370",X"00ED",X"FE1D",X"FDF1",X"FEAD",X"FED8",X"FF26",X"FF0F",X"FE39",X"FE09",X"FE29",X"FE43",X"FF02",X"0155",X"034F",X"0452",X"0426",X"02C0",X"FF9E",X"FDE1",X"FE61",X"FEC4",X"FF08",X"FF74",X"FEB5",X"FE19",X"FE1B",X"FE39",X"FE4A",X"FFC4",X"020D",X"03BB",X"0451",X"0412",X"01CA",X"FEC6",X"FE15",X"FE99",X"FEB5",X"FF43",X"FF2F",X"FE66",X"FE11",X"FE39",X"FE13",X"FE94",X"008D",X"02B4",X"040A",X"046F",X"039D",X"007E",X"FE55",X"FE51",X"FE94",X"FEEF",X"FF59",X"FEC1",X"FE22",X"FE0C",X"FE2F",X"FDFB",X"FF1C",X"013D",X"0336",X"042D",X"0495",X"02AA",X"FF85",X"FE68",X"FEA0",X"FEAE",X"FF53",X"FF46",X"FE92",X"FE05",X"FE3D",X"FDFB",X"FE35",X"FFBC",X"01FE",X"0363",X"046B",X"0419",X"0152",X"FED1",X"FE7E",X"FE77",X"FEDD",X"FF67",X"FF15",X"FE4C",X"FE3B",X"FE3E",X"FE06",X"FEB5",X"00B7",X"0292",X"03D4",X"04C2",X"0344",X"0022",X"FE9E",X"FE65",X"FE82",X"FF1A",X"FF59",X"FEB4",X"FE2B",X"FE49",X"FE0E",X"FE19",X"FF4A",X"0168",X"02E4",X"045C",X"049C",X"0210",X"FF77",X"FEA6",X"FE62",X"FED3",X"FF5E",X"FF36",X"FE54",X"FE41",X"FE2A",X"FDF0",X"FE42",X"001E",X"01DC",X"0347",X"04C6",X"03FB",X"00F8",X"FF2F",X"FE81",X"FE82",X"FF16",X"FF83",X"FED3",X"FE3D",X"FE3A",X"FE17",X"FDD3",X"FEDB",X"00BA",X"022F",X"03F7",X"04D3",X"02C1",X"0027",X"FEEF",X"FE74",X"FEA8",X"FF76",X"FF5C",X"FE80",X"FE3E",X"FE2D",X"FDE6",X"FE00",X"FF9A",X"012E",X"02B4",X"04A8",X"047A",X"01D4",X"FFC0",X"FEAD",X"FE79",X"FEFD",X"FF96",X"FF00",X"FE5E",X"FE3A",X"FE2B",X"FDAA",X"FE7F",X"0029",X"0192",X"0387",X"050D",X"037B",X"010F",X"FF4D",X"FE80",X"FE7E",X"FF59",X"FF65",X"FEA4",X"FE31",X"FE4C",X"FDDA",X"FDCA",X"FF26",X"009A",X"0217",X"046E",X"04AB",X"0293",X"0058",X"FF0B",X"FE73",X"FEF5",X"FF8F",X"FF2F",X"FE74",X"FE49",X"FE3D",X"FDA7",X"FE30",X"FF9D",X"00C6",X"02E3",X"04CA",X"0405",X"01BF",X"FFE0",X"FEBB",X"FE7B",X"FF4D",X"FF77",X"FECD",X"FE3A",X"FE59",X"FDEF",X"FDBB",X"FEDF",X"FFEB",X"015D",X"03DF",X"04CE",X"034D",X"0112",X"FF8F",X"FE81",X"FEE3",X"FF82",X"FF56",X"FE70",X"FE50",X"FE35",X"FDA3",X"FDF7",X"FF36",X"0006",X"0235",X"047D",X"047B",X"027F",X"00A1",X"FF17",X"FE9B",X"FF33",X"FF9B",X"FEF4",X"FE57",X"FE61",X"FDEE",X"FD84",X"FE8B",X"FF55",X"00AC",X"033B",X"04CE",X"03C6",X"01C3",X"FFF6",X"FEB2",X"FEC1",X"FF7B",X"FF86",X"FEAF",X"FE74",X"FE5B",X"FD90",X"FDE4",X"FEEA",X"FF96",X"0189",X"0409",X"04A6",X"030C",X"0124",X"FF59",X"FE96",X"FF07",X"FFB5",X"FF31",X"FE91",X"FE92",X"FE0E",X"FD7A",X"FE5F",X"FEDE",X"0001",X"0277",X"0488",X"041B",X"027C",X"0084",X"FEF2",X"FEA5",X"FF67",X"FFA6",X"FEE0",X"FE8D",X"FE81",X"FD87",X"FDB6",X"FE75",X"FF09",X"00C6",X"0396",X"04AE",X"03B3",X"01ED",X"FFE5",X"FEA9",X"FEF6",X"FFBE",X"FF5E",X"FE9A",X"FEA8",X"FDF0",X"FD60",X"FE04",X"FE94",X"FF5B",X"01CA",X"0434",X"0473",X"032A",X"0129",X"FF63",X"FEA6",X"FF61",X"FFC3",X"FEF5",X"FEBA",X"FE95",X"FDA1",X"FDBE",X"FE4D",X"FE9F",X"FFF7",X"02D4",X"0460",X"0408",X"027E",X"006E",X"FED8",X"FED4",X"FFB6",X"FF82",X"FEC8",X"FEEC",X"FE1C",X"FD8C",X"FDFF",X"FE6C",X"FED7",X"00FF",X"0389",X"047B",X"0391",X"01C3",X"FFAD",X"FE9E",X"FF37",X"FFDE",X"FF19",X"FEFD",X"FEB3",X"FDC3",X"FDA6",X"FE2C",X"FE48",X"FF5A",X"0202",X"0419",X"0457",X"0322",X"0112",X"FF34",X"FED4",X"FFBF",X"FFAD",X"FF10",X"FF11",X"FE3E",X"FD8D",X"FDDE",X"FE2A",X"FE3C",X"0028",X"02BF",X"043A",X"03F1",X"0270",X"004D",X"FED8",X"FF41",X"FFF6",X"FF53",X"FF47",X"FEEE",X"FDF9",X"FDA4",X"FE29",X"FDFB",X"FECE",X"011C",X"0366",X"0432",X"0387",X"01B6",X"FFA0",X"FECD",X"FFBC",X"FFAA",X"FF44",X"FF3C",X"FE83",X"FDA4",X"FDF3",X"FE1E",X"FDFA",X"FF6A",X"01FB",X"03D6",X"042E",X"031C",X"010C",X"FF0F",X"FF3F",X"FFCC",X"FF62",X"FF51",X"FF0B",X"FE03",X"FDB4",X"FE1B",X"FDD4",X"FE39",X"0038",X"02B7",X"0417",X"0402",X"0296",X"0041",X"FF12",X"FFBB",X"FF9C",X"FF64",X"FF6A",X"FEB5",X"FDB8",X"FDF3",X"FE02",X"FDB8",X"FEAD",X"0116",X"033D",X"041E",X"0399",X"01B5",X"FF66",X"FF56",X"FFB9",X"FF75",X"FF8A",X"FF68",X"FE53",X"FDF3",X"FE3D",X"FDF4",X"FDF0",X"FF7F",X"01E6",X"03A2",X"0406",X"0325",X"00AC",X"FF44",X"FF8E",X"FF9B",X"FF6A",X"FF91",X"FEEC",X"FDF8",X"FE17",X"FE31",X"FDC8",X"FE55",X"005F",X"02C2",X"03EE",X"0413",X"0258",X"FFE2",X"FF4A",X"FFA2",X"FF6F",X"FF76",X"FF6C",X"FE6A",X"FDEC",X"FE2E",X"FDE9",X"FDAA",X"FEE0",X"0138",X"032D",X"042E",X"03D0",X"015A",X"FFB1",X"FFA3",X"FFA8",X"FF76",X"FFC1",X"FF18",X"FE14",X"FE08",X"FE15",X"FDA1",X"FDD5",X"FF8A",X"01EA",X"038A",X"0462",X"02F5",X"0072",X"FF8E",X"FFB0",X"FF80",X"FFB1",X"FFBC",X"FEA9",X"FE00",X"FE33",X"FDE9",X"FD8C",X"FE44",X"0076",X"026E",X"0404",X"0425",X"01FC",X"0000",X"FFC4",X"FFA9",X"FF86",X"FFE0",X"FF4F",X"FE3D",X"FE0B",X"FE1F",X"FDB4",X"FD98",X"FF08",X"0124",X"0301",X"046F",X"0376",X"0118",X"FFF1",X"FFCA",X"FF8D",X"FFC1",X"FFD6",X"FEDB",X"FE14",X"FE22",X"FE00",X"FD85",X"FDE1",X"FFD2",X"01A1",X"03B9",X"0465",X"029B",X"007C",X"FFFF",X"FFA9",X"FF95",X"FFF8",X"FF94",X"FE6A",X"FE28",X"FE2B",X"FDCC",X"FD53",X"FE8C",X"004F",X"0246",X"0435",X"03DE",X"0193",X"003E",X"FFEC",X"FF97",X"FFD4",X"000D",X"FF12",X"FE3B",X"FE35",X"FE29",X"FD70",X"FD9D",X"FF29",X"00DF",X"0329",X"0482",X"032A",X"0113",X"003D",X"FFB9",X"FF92",X"0006",X"FFB1",X"FE9F",X"FE2C",X"FE57",X"FDF8",X"FD5A",X"FE34",X"FF98",X"018A",X"03D6",X"0437",X"0235",X"00B3",X"001A",X"FF93",X"FFD0",X"0033",X"FF50",X"FE62",X"FE39",X"FE46",X"FD79",X"FD87",X"FE9E",X"001E",X"0273",X"0465",X"0377",X"018F",X"0087",X"FFE7",X"FF99",X"002C",X"FFEE",X"FEEC",X"FE2D",X"FE6B",X"FDF4",X"FD5C",X"FDE1",X"FF04",X"00C5",X"036C",X"0448",X"02B1",X"0129",X"004F",X"FF9A",X"FFD4",X"002F",X"FF98",X"FE85",X"FE4C",X"FE5B",X"FD94",X"FD87",X"FE47",X"FF87",X"01D2",X"0421",X"03D7",X"021D",X"00E6",X"0001",X"FF98",X"0011",X"0012",X"FF2D",X"FE44",X"FE71",X"FDF9",X"FD6C",X"FDBA",X"FE88",X"000F",X"02D9",X"043C",X"032D",X"019B",X"0098",X"FFA9",X"FFDF",X"0040",X"FFEB",X"FEB6",X"FE65",X"FE5A",X"FDAA",X"FD70",X"FE04",X"FECE",X"0109",X"03A0",X"03FE",X"0278",X"0166",X"002B",X"FFBE",X"0026",X"0065",X"FF71",X"FE81",X"FE8B",X"FE22",X"FD76",X"FDA6",X"FE26",X"FF5A",X"0213",X"0406",X"0360",X"0210",X"00D2",X"FFDA",X"FFC5",X"0057",X"0038",X"FEF4",X"FE8E",X"FE7D",X"FDCA",X"FD83",X"FDCA",X"FE40",X"0038",X"030B",X"03F1",X"02ED",X"01C0",X"0065",X"FFC2",X"0004",X"0091",X"FFB6",X"FEC3",X"FEB2",X"FE41",X"FD86",X"FDA4",X"FDC9",X"FEA9",X"014F",X"03A6",X"03A1",X"02A3",X"0139",X"001C",X"FFB9",X"006B",X"007E",X"FF43",X"FEBA",X"FE91",X"FDD4",X"FD7B",X"FDA2",X"FDCD",X"FF54",X"024A",X"03A3",X"0347",X"0223",X"00CE",X"FFD3",X"FFF9",X"00BD",X"0016",X"FF18",X"FEF1",X"FE7D",X"FDC9",X"FDC0",X"FDAA",X"FE10",X"0078",X"030B",X"03A1",X"02F4",X"01A4",X"004D",X"FFAF",X"0069",X"008E",X"FF85",X"FEF3",X"FEC9",X"FDFF",X"FDA0",X"FD99",X"FD78",X"FEA0",X"01A1",X"035F",X"0394",X"028E",X"0147",X"FFE6",X"FFE5",X"00AD",X"0046",X"FF47",X"FF1A",X"FE9B",X"FDE3",X"FDC8",X"FD9C",X"FD8F",X"FFAC",X"0253",X"0387",X"0342",X"0230",X"00AB",X"FFB1",X"004C",X"00B6",X"FFB9",X"FF2A",X"FEFA",X"FE3E",X"FDCE",X"FDCF",X"FD5A",X"FE20",X"00BA",X"02D4",X"037D",X"02E3",X"01A3",X"0014",X"FFCE",X"009E",X"005D",X"FF75",X"FF46",X"FEC3",X"FE0A",X"FE05",X"FDAC",X"FD5A",X"FEFE",X"0187",X"0341",X"0370",X"02AA",X"0113",X"FFD6",X"0032",X"00BD",X"FFE8",X"FF69",X"FF1A",X"FE59",X"FDE3",X"FDF1",X"FD36",X"FDB5",X"FFE3",X"024A",X"0354",X"033F",X"0231",X"007A",X"FFDE",X"00B0",X"0083",X"FFB2",X"FF67",X"FEDB",X"FDFD",X"FE04",X"FD9A",X"FD18",X"FE46",X"00CB",X"02D9",X"0372",X"031E",X"019A",X"FFFC",X"0041",X"00D0",X"0028",X"FF9B",X"FF60",X"FE72",X"FE06",X"FE00",X"FD37",X"FD4A",X"FF12",X"019C",X"030A",X"0367",X"02A7",X"00D3",X"FFF7",X"00A9",X"009F",X"FFE3",X"FF99",X"FF1A",X"FE27",X"FE2B",X"FDBB",X"FD15",X"FDD4",X"0015",X"0241",X"0358",X"0362",X"020A",X"003C",X"003E",X"00B6",X"004A",X"FFC8",X"FF97",X"FE9A",X"FE28",X"FE19",X"FD61",X"FD11",X"FE84",X"00E9",X"02AE",X"0373",X"031E",X"012D",X"001A",X"007F",X"00AB",X"0000",X"FFF3",X"FF50",X"FE66",X"FE5A",X"FDE5",X"FD11",X"FD4F",X"FF51",X"017D",X"02E3",X"0384",X"0265",X"008D",X"0050",X"00DC",X"0086",X"0019",X"FFE9",X"FEEA",X"FE77",X"FE52",X"FD92",X"FCDD",X"FDDB",X"FFFB",X"01E3",X"0333",X"034C",X"0187",X"0033",X"0091",X"00BC",X"0033",X"002D",X"FF8D",X"FEB1",X"FE91",X"FE33",X"FD37",X"FD18",X"FE96",X"00B2",X"0264",X"0397",X"02D3",X"00EB",X"0049",X"00CB",X"007C",X"003B",X"0005",X"FF25",X"FE92",X"FE7E",X"FDC7",X"FCE8",X"FD6E",X"FF5E",X"013E",X"02FF",X"039B",X"0224",X"0079",X"00AB",X"00C0",X"005B",X"0061",X"FFAC",X"FEC3",X"FE8F",X"FE4C",X"FD5F",X"FCD4",X"FE11",X"FFFA",X"01D5",X"0379",X"0337",X"0149",X"0086",X"00DB",X"007D",X"0076",X"0030",X"FF5C",X"FEB4",X"FEAD",X"FE1F",X"FD14",X"FD2A",X"FEBA",X"006D",X"0277",X"0395",X"0270",X"00A9",X"00AE",X"009E",X"0075",X"007C",X"FFE9",X"FF03",X"FECC",X"FEA1",X"FDBC",X"FCD7",X"FDB5",X"FF3E",X"012C",X"0327",X"0380",X"01A0",X"00B3",X"00C6",X"0089",X"0086",X"005F",X"FF82",X"FEDB",X"FEC5",X"FE5F",X"FD3B",X"FD13",X"FE3F",X"FFBD",X"01EC",X"0394",X"02C6",X"010C",X"00D2",X"00A6",X"0079",X"0090",X"0024",X"FF34",X"FED4",X"FECA",X"FDF5",X"FCF4",X"FD73",X"FEA0",X"0058",X"02A7",X"038D",X"01FF",X"00F9",X"00E2",X"00A5",X"00AD",X"0099",X"FFD1",X"FF1A",X"FEFA",X"FEA6",X"FD60",X"FD00",X"FDBF",X"FF17",X"0132",X"0357",X"02F5",X"0164",X"00D8",X"00A1",X"0082",X"00AB",X"004E",X"FF74",X"FEF8",X"FF0C",X"FE38",X"FD2D",X"FD51",X"FE3B",X"FFA9",X"0233",X"0387",X"0252",X"013E",X"00E0",X"0092",X"00AD",X"00BA",X"0008",X"FF1A",X"FEFF",X"FEBE",X"FDA3",X"FD17",X"FD91",X"FE79",X"0072",X"030A",X"0327",X"01C9",X"011A",X"00C3",X"00A1",X"00D5",X"0099",X"FFAF",X"FF00",X"FF0D",X"FE53",X"FD68",X"FD37",X"FDCC",X"FEF9",X"0193",X"0353",X"0293",X"0183",X"00FB",X"00AA",X"00C4",X"00E4",X"0066",X"FF59",X"FF2F",X"FEF5",X"FDEB",X"FD31",X"FD64",X"FDE1",X"FFC5",X"0276",X"0320",X"0215",X"013F",X"00B9",X"009C",X"00D6",X"00EE",X"FFF1",X"FF3D",X"FF49",X"FEA7",X"FD94",X"FD48",X"FD7C",X"FE47",X"00E1",X"02FD",X"02C5",X"01CD",X"0102",X"009F",X"00A4",X"00F8",X"0097",X"FF98",X"FF59",X"FF2D",X"FE35",X"FD65",X"FD78",X"FD79",X"FF16",X"01DF",X"030E",X"026A",X"0192",X"00E3",X"00A0",X"00CC",X"0105",X"0024",X"FF80",X"FF63",X"FEDE",X"FDB1",X"FD6B",X"FD47",X"FDB3",X"0016",X"027F",X"02DE",X"021E",X"014A",X"00C8",X"00AE",X"010F",X"00BE",X"FFCB",X"FF73",X"FF5F",X"FE5C",X"FD83",X"FD68",X"FD35",X"FE6C",X"0136",X"02D5",X"02A0",X"01C7",X"010C",X"0095",X"00CF",X"011D",X"005F",X"FF9C",X"FF93",X"FF12",X"FDFE",X"FDAC",X"FD4A",X"FD4C",X"FF67",X"01F2",X"02C5",X"0248",X"0180",X"00C8",X"0090",X"010C",X"00ED",X"FFFF",X"FF8F",X"FF89",X"FE96",X"FDDC",X"FDAF",X"FD1A",X"FDD8",X"007E",X"0272",X"02C3",X"0217",X"0150",X"0087",X"00B9",X"011D",X"0095",X"FFB4",X"FFB4",X"FF3D",X"FE2B",X"FDC8",X"FD5C",X"FCFA",X"FEC7",X"0143",X"02A9",X"027A",X"01DF",X"00F7",X"0097",X"0116",X"012A",X"0041",X"FFD1",X"FFCC",X"FED6",X"FE0A",X"FDD6",X"FCF0",X"FD4F",X"FF9C",X"01E0",X"029C",X"0237",X"016C",X"009B",X"00AC",X"0136",X"00C2",X"FFF9",X"FFF1",X"FF78",X"FE77",X"FE2C",X"FD8F",X"FCD4",X"FE1B",X"008B",X"0251",X"0281",X"020D",X"010C",X"008F",X"00FD",X"012B",X"0057",X"FFF1",X"FFE3",X"FF05",X"FE51",X"FE1D",X"FD24",X"FD1B",X"FEF0",X"0150",X"025A",X"0263",X"01AB",X"00C2",X"00A4",X"012C",X"00DB",X"0020",X"0014",X"FFA5",X"FE9D",X"FE74",X"FDBF",X"FCDD",X"FD7A",X"FFC4",X"01B9",X"026A",X"0234",X"0145",X"0086",X"00DF",X"013E",X"0087",X"0028",X"0038",X"FF44",X"FEAC",X"FE6B",X"FD54",X"FCD0",X"FE31",X"009A",X"0204",X"0275",X"01F0",X"00E8",X"0092",X"0131",X"010A",X"0040",X"004D",X"FFE4",X"FEE3",X"FEA7",X"FE05",X"FCF9",X"FD10",X"FF28",X"013B",X"0254",X"0268",X"0199",X"0099",X"00D8",X"0134",X"008E",X"0034",X"0048",X"FF6A",X"FEE3",X"FE97",X"FDA3",X"FCB3",X"FDBB",X"FFF6",X"01AF",X"027E",X"0243",X"0110",X"008C",X"011D",X"00FE",X"0053",X"007B",X"FFFC",X"FF22",X"FEE4",X"FE69",X"FD25",X"FCD3",X"FE7E",X"0095",X"0200",X"0281",X"01CF",X"00B2",X"00D1",X"0153",X"00B0",X"0069",X"007A",X"FF9E",X"FF11",X"FEE4",X"FDE1",X"FCC3",X"FD3D",X"FF37",X"0124",X"024B",X"0270",X"0143",X"008B",X"0120",X"0116",X"007F",X"00AA",X"0033",X"FF6B",X"FF09",X"FEB9",X"FD61",X"FCB5",X"FDD7",X"FFEA",X"0196",X"0282",X"0206",X"00CF",X"00BC",X"0145",X"00BF",X"009A",X"008C",X"FFD8",X"FF31",X"FF29",X"FE56",X"FCFB",X"FD03",X"FE9E",X"0082",X"01FB",X"0272",X"0183",X"00A9",X"0121",X"0122",X"00A3",X"00C0",X"0062",X"FF88",X"FF40",X"FEFA",X"FDB6",X"FCB1",X"FD66",X"FF40",X"0101",X"0255",X"023C",X"0100",X"00CD",X"0142",X"00C7",X"00C7",X"00B8",X"000A",X"FF5F",X"FF50",X"FE9A",X"FD38",X"FCD5",X"FE13",X"FFD8",X"019A",X"0271",X"01A5",X"00B7",X"012B",X"010F",X"00C3",X"00E5",X"009D",X"FFBF",X"FF61",X"FF35",X"FE10",X"FCDC",X"FD2A",X"FEA6",X"0068",X"0216",X"0251",X"011D",X"00EF",X"0133",X"00EB",X"00CA",X"00ED",X"0041",X"FF7D",X"FF5E",X"FEDE",X"FD7A",X"FCCA",X"FDA5",X"FF4A",X"011C",X"0278",X"01E6",X"00F6",X"012C",X"010F",X"00B6",X"00D8",X"00B2",X"FFD5",X"FF70",X"FF74",X"FE7D",X"FD23",X"FD04",X"FE26",X"FFD9",X"01BF",X"0269",X"013F",X"00F4",X"0122",X"00D5",X"00CA",X"0100",X"007F",X"FFA7",X"FF9F",X"FF50",X"FDEC",X"FCF8",X"FD49",X"FE9B",X"0079",X"0235",X"01E1",X"011A",X"0126",X"010E",X"00B6",X"00F6",X"00E8",X"0021",X"FF94",X"FFA6",X"FED5",X"FD6F",X"FCF9",X"FDB3",X"FF28",X"0156",X"0240",X"0173",X"011E",X"0134",X"00DD",X"00C5",X"0119",X"0097",X"FFD6",X"FFB7",X"FF8E",X"FE4D",X"FD1A",X"FD23",X"FDFD",X"FFDB",X"01EA",X"01E9",X"012D",X"0122",X"0104",X"00B1",X"00F9",X"0103",X"0053",X"FFD0",X"FFEC",X"FF46",X"FDDA",X"FD1B",X"FD61",X"FE7B",X"00D3",X"0211",X"0185",X"0118",X"0123",X"00D6",X"00C4",X"0117",X"00D2",X"FFFD",X"FFDC",X"FFC7",X"FEB6",X"FD67",X"FD27",X"FD7F",X"FF54",X"0187",X"01EE",X"0148",X"0139",X"0117",X"00B0",X"00F5",X"0124",X"007C",X"FFE1",X"FFE5",X"FF8C",X"FE1E",X"FD3E",X"FD1B",X"FDF2",X"003B",X"01DA",X"019E",X"0124",X"0135",X"00DD",X"00BB",X"0130",X"010A",X"0039",X"FFF2",X"FFF7",X"FF1A",X"FDC3",X"FD2F",X"FD18",X"FEA5",X"00FB",X"01C2",X"0148",X"0141",X"010D",X"00BC",X"00E3",X"0158",X"00C9",X"0018",X"0014",X"FFDA",X"FE70",X"FD92",X"FD0E",X"FD75",X"FF9F",X"0179",X"0185",X"013F",X"0139",X"00E9",X"00A4",X"0135",X"013A",X"0076",X"0015",X"003E",X"FF57",X"FE19",X"FD63",X"FCF0",X"FE2B",X"0074",X"0183",X"014C",X"0139",X"010E",X"0092",X"00DA",X"014F",X"0103",X"0030",X"0035",X"000C",X"FEDD",X"FDE6",X"FD16",X"FD37",X"FF11",X"010F",X"0173",X"014E",X"0142",X"00D6",X"0093",X"011E",X"0157",X"00A5",X"0029",X"0056",X"FFA1",X"FE98",X"FD94",X"FCDE",X"FDA1",X"FFDE",X"0139",X"0148",X"0149",X"0129",X"0090",X"00B3",X"0152",X"0121",X"0058",X"0067",X"003A",X"FF4E",X"FE6A",X"FD5E",X"FCEE",X"FE82",X"0089",X"0140",X"013B",X"0150",X"00DF",X"0072",X"00DA",X"014D",X"00BB",X"004A",X"007F",X"FFD9",X"FEFF",X"FE0A",X"FCEC",X"FD5F",X"FF70",X"00F8",X"0136",X"0160",X"013A",X"00A3",X"008F",X"0140",X"013A",X"006C",X"0073",X"0044",X"FF81",X"FEB5",X"FD79",X"FCB0",X"FE05",X"000D",X"0114",X"0154",X"0178",X"010B",X"008B",X"00D6",X"0169",X"00E9",X"0069",X"0081",X"FFFE",X"FF4C",X"FE62",X"FCFC",X"FD04",X"FECD",X"0086",X"0101",X"015A",X"0157",X"00B9",X"0078",X"012E",X"014B",X"00A1",X"009B",X"0067",X"FFCD",X"FF25",X"FDDB",X"FCC0",X"FD87",X"FF98",X"00C0",X"0123",X"016F",X"0128",X"007E",X"00B0",X"0156",X"00EC",X"008B",X"00A5",X"0024",X"FFA7",X"FEBC",X"FD3F",X"FCC6",X"FE56",X"001A",X"00E5",X"015A",X"0170",X"00DA",X"005D",X"0108",X"0144",X"00AB",X"0096",X"006D",X"FFF5",X"FF79",X"FE37",X"FCD5",X"FD43",X"FF1E",X"006A",X"0119",X"0189",X"0160",X"0090",X"0097",X"012C",X"00F5",X"00A7",X"009C",X"003A",X"FFEC",X"FF31",X"FDA3",X"FCAE",X"FDE4",X"FF91",X"008A",X"012E",X"018C",X"00ED",X"0055",X"00F2",X"0143",X"00D7",X"00CE",X"0094",X"0035",X"FFE6",X"FEBF",X"FD0E",X"FCF5",X"FE94",X"FFEF",X"00BD",X"015B",X"0164",X"0084",X"007B",X"011B",X"00FF",X"00D6",X"00C9",X"006C",X"0033",X"FFB2",X"FE0D",X"FCC8",X"FD83",X"FF15",X"002C",X"00E7",X"0186",X"0106",X"0050",X"00C9",X"0122",X"00D9",X"00DF",X"009D",X"005E",X"003D",X"FF46",X"FD61",X"FCD7",X"FE11",X"FF85",X"0072",X"0152",X"0184",X"009A",X"006E",X"010B",X"00FC",X"00E3",X"00D4",X"006C",X"0052",X"001A",X"FE92",X"FCF4",X"FD3D",X"FEB4",X"FFC1",X"00A1",X"017B",X"011E",X"0064",X"00AC",X"0102",X"00F4",X"00FF",X"00A8",X"0067",X"0079",X"FFBE");
begin
 
   
 process(resetN, CLK)
	 type noteArrd is array (0 to 12) of integer;
	 variable dataTmp : noteArrd;
 begin
	if (resetN='0') then
		dataTmp := (others  => 0);
	elsif(rising_edge(CLK)) then
		dataTmp := (others  => 0);
		for i in 0 to 12 loop
			if conv_integer(addrArr(i)) > 0 then
				dataTmp(i) := conv_integer(sound0(conv_integer(addrArr(i))));
			end if;
		end loop;
	end if;
	Q <= conv_std_logic_vector(dataTmp(0) + dataTmp(1) + dataTmp(2) + dataTmp(3) + dataTmp(4) + dataTmp(5) + dataTmp(6) + dataTmp(7) + dataTmp(8) + dataTmp(9) + dataTmp(10) + dataTmp(11) + dataTmp(12), 16);
end process;
	 

		   
end arch;