--------------------------------------
-- SinTable.vhd
-- Written by Gadi and Eran Tuchman.
-- All rights reserved, Copyright 2009
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all ;

entity sintable is
port(
  CLK     					: in std_logic;
  resetN 					: in std_logic;
  ADDR    					: in std_logic_vector(13 downto 0);
  Q       					: out std_logic_vector(15 downto 0)
);
end sintable;

architecture arch of sintable is
constant array_size 			: integer := 14700 ;

type table_type is array(0 to array_size - 1) of std_logic_vector(15 downto 0);
signal sin_table				: table_type;
signal Q_tmp       			:  std_logic_vector(15 downto 0) ;



begin
 
   
  sintable_proc: process(resetN, CLK)
    constant sin_table : table_type := (X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"FFFF",X"0000",X"0000",X"0000",X"0000",X"FFFF",X"0000",X"0000",X"0000",X"FFFF",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"FFFF",X"FFFF",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"FFFE",X"0000",X"0000",X"0000",X"0000",X"FFFF",X"0000",X"0000",X"0000",X"0000",X"FFFF",X"FFFD",X"FFFD",X"0000",X"0001",X"0000",X"0000",X"0000",X"FFFF",X"FFFF",X"FFFF",X"FFFE",X"FFFE",X"FFFD",X"FFFE",X"0000",X"0007",X"0006",X"0006",X"FFFF",X"0004",X"FFFE",X"0000",X"FFF5",X"FFFE",X"FFF3",X"0002",X"0004",X"0004",X"FFF3",X"FFF9",X"FFFD",X"0005",X"0012",X"0005",X"0013",X"000C",X"FFFA",X"0002",X"FFFF",X"FFFE",X"FFFC",X"FFFB",X"FFFC",X"FFFB",X"0006",X"FFF9",X"FFF9",X"FFFD",X"0005",X"0004",X"0000",X"0001",X"0002",X"0007",X"FFF8",X"FFF9",X"FFF4",X"0003",X"0002",X"FFF6",X"FFF9",X"0000",X"0012",X"0006",X"FFFF",X"0002",X"0000",X"0003",X"0003",X"FFFE",X"0003",X"0000",X"000E",X"0005",X"FFFD",X"0001",X"FFFB",X"FFFC",X"0000",X"FFFA",X"0006",X"FFF8",X"0002",X"FFFE",X"FFFA",X"0004",X"0000",X"0003",X"0000",X"0000",X"FFF8",X"0000",X"0001",X"FFFF",X"FFF9",X"0003",X"FFFA",X"FFF5",X"FFFE",X"FFFD",X"FFFD",X"0001",X"000E",X"0000",X"0004",X"0008",X"000E",X"000A",X"0000",X"0003",X"FFFE",X"FFFB",X"FFFC",X"FFFE",X"FFFF",X"0009",X"0001",X"FFFF",X"0009",X"FFFF",X"0000",X"FFF6",X"0001",X"FFFF",X"FFF9",X"FFFC",X"FFFF",X"FFFB",X"0000",X"FFFA",X"FFF1",X"FFFC",X"FFFC",X"FFF4",X"0001",X"0004",X"0008",X"0006",X"0008",X"0005",X"0001",X"000C",X"0008",X"0001",X"0009",X"0000",X"FFF5",X"0008",X"0008",X"FFFE",X"FFFF",X"0001",X"FFF9",X"FFFD",X"FFFD",X"FFF0",X"FFF9",X"FFF7",X"0000",X"FFFB",X"FFFC",X"0001",X"0002",X"000A",X"FFFB",X"0005",X"0004",X"0000",X"0000",X"0005",X"0001",X"0001",X"000E",X"FFFE",X"FFF3",X"FFF6",X"FFFF",X"FFEE",X"FFF9",X"FFFC",X"FFFD",X"FFFC",X"FFFA",X"0008",X"000A",X"000D",X"0008",X"0002",X"0007",X"000A",X"0004",X"FFFE",X"FFFD",X"FFFC",X"FFFC",X"FFF2",X"0000",X"FFFE",X"0005",X"FFFF",X"0006",X"000D",X"0006",X"FFF9",X"000B",X"FFFF",X"FFF8",X"0004",X"FFFC",X"FFF5",X"0003",X"FFF6",X"0000",X"0003",X"FFFC",X"0003",X"FFF6",X"FFF6",X"FFF9",X"FFFF",X"FFF8",X"FFF6",X"0001",X"FFFF",X"0000",X"FFFD",X"0005",X"000C",X"0007",X"000D",X"000A",X"FFFF",X"FFF8",X"0004",X"0005",X"FFFF",X"FFFE",X"FFFB",X"FFFC",X"FFF7",X"FFFE",X"0004",X"FFFF",X"FFF9",X"0001",X"0000",X"0000",X"FFFF",X"0000",X"FFFC",X"FFFA",X"FFFF",X"FFF8",X"000B",X"FFFF",X"FFFC",X"FFF9",X"0004",X"FFFD",X"0008",X"FFFD",X"FFFC",X"FFF5",X"0006",X"0000",X"0003",X"0007",X"0000",X"0007",X"0003",X"0000",X"FFF7",X"FFFF",X"FFF6",X"FFFC",X"0005",X"0000",X"FFFC",X"0000",X"FFF4",X"0000",X"FFF7",X"FFFD",X"FFFE",X"0000",X"0009",X"0004",X"0005",X"FFFF",X"FFFF",X"FFFD",X"0000",X"FFFE",X"FFFE",X"0001",X"0001",X"FFF5",X"FFFA",X"FFF9",X"FFF8",X"0000",X"FFFB",X"FFF7",X"0000",X"0003",X"0007",X"0001",X"0000",X"000F",X"0003",X"0004",X"0009",X"FFFE",X"FFFF",X"FFFA",X"FFFC",X"FFFC",X"0004",X"0003",X"FFFC",X"FFFC",X"FFFC",X"FFFA",X"0006",X"FFF2",X"FFF9",X"0003",X"FFFF",X"FFFF",X"0002",X"0004",X"0001",X"0003",X"0002",X"FFF8",X"FFFE",X"FFFB",X"FFF8",X"0001",X"0001",X"0004",X"FFFF",X"FFFE",X"FFFE",X"0002",X"000B",X"0000",X"FFFB",X"FFFC",X"FFF7",X"FFF8",X"FFFC",X"FFFA",X"FFFC",X"0000",X"0002",X"0007",X"FFF8",X"FFF9",X"FFFA",X"FFFF",X"0002",X"0009",X"FFFF",X"0004",X"FFF7",X"FFFE",X"FFFF",X"0001",X"FFFC",X"FFFE",X"0007",X"0001",X"0001",X"0002",X"FFFA",X"0006",X"0002",X"FFFE",X"FFFC",X"0006",X"0007",X"0000",X"0002",X"0006",X"FFF5",X"0002",X"FFFC",X"0002",X"0007",X"0000",X"0015",X"FFFE",X"FFFC",X"0004",X"0007",X"0005",X"0007",X"0006",X"FFF0",X"FFF9",X"FFFD",X"FFFD",X"FFF8",X"FFFE",X"FFF4",X"FFFF",X"FFFF",X"0014",X"000A",X"0002",X"0004",X"0008",X"FFFF",X"0007",X"0005",X"0004",X"FFFA",X"0005",X"FFFA",X"0003",X"FFF8",X"FFF8",X"FFFC",X"0000",X"FFF6",X"FFFD",X"0002",X"0005",X"FFFB",X"FFFE",X"0000",X"0000",X"0000",X"FFFD",X"FFFD",X"0003",X"FFFA",X"0004",X"0009",X"0008",X"FFFD",X"0001",X"FFFF",X"0002",X"FFF7",X"FFFB",X"FFEE",X"FFF3",X"FFFE",X"FFF9",X"0000",X"0004",X"0005",X"0003",X"0002",X"0001",X"0005",X"FFFD",X"0004",X"FFFD",X"0000",X"FFFF",X"FFFD",X"FFFF",X"FFFC",X"FFFB",X"FFF7",X"0001",X"FFF2",X"FFFA",X"FFFC",X"0003",X"0002",X"0004",X"0007",X"0005",X"0008",X"FFFE",X"0002",X"0001",X"FFF5",X"FFF6",X"0001",X"0005",X"0006",X"FFFC",X"FFFF",X"0000",X"FFF9",X"FFFD",X"FFFC",X"0000",X"0002",X"FFF7",X"FFF8",X"FFFF",X"FFFA",X"FFFE",X"0000",X"FFFD",X"0000",X"FFFF",X"0002",X"FFFA",X"0000",X"FFFA",X"0006",X"0004",X"0004",X"000C",X"0004",X"0008",X"0003",X"FFFE",X"FFFE",X"0002",X"FFFC",X"0003",X"FFFB",X"FFFD",X"0001",X"0004",X"FFF7",X"FFF1",X"FFFF",X"FFFD",X"0004",X"0000",X"FFFD",X"FFFE",X"0000",X"0000",X"FFFE",X"0005",X"0000",X"0000",X"0001",X"0003",X"0007",X"000B",X"FFFD",X"0000",X"0001",X"FFFE",X"FFFE",X"0001",X"FFFB",X"0000",X"0005",X"FFF9",X"FFF6",X"0001",X"FFFE",X"FFF8",X"FFF4",X"FFFF",X"FFFC",X"FFF8",X"FFFD",X"000C",X"0008",X"FFFD",X"FFFC",X"0003",X"0007",X"0000",X"000D",X"0009",X"0004",X"0001",X"0001",X"FFFE",X"FFFD",X"FFED",X"FFFD",X"FFFE",X"0005",X"FFFC",X"0007",X"000C",X"FFFC",X"0009",X"0007",X"0006",X"0004",X"0000",X"FFFD",X"0000",X"FFFC",X"0007",X"FFFB",X"0000",X"FFF9",X"FFFC",X"FFF7",X"FFFC",X"FFFD",X"FFF6",X"0004",X"FFFC",X"0003",X"0001",X"0000",X"000B",X"000F",X"FFFF",X"FFFE",X"FFF7",X"000B",X"FFFE",X"FFFB",X"FFFC",X"FFEF",X"FFFA",X"0000",X"FFFF",X"0002",X"FFFB",X"FFFE",X"0000",X"FFF6",X"FFFF",X"000C",X"0002",X"0003",X"0006",X"FFFF",X"FFFE",X"000A",X"0006",X"0007",X"0007",X"FFFD",X"FFFD",X"FFFC",X"FFEF",X"FFF2",X"FFF8",X"0000",X"0000",X"FFFB",X"0000",X"FFFE",X"000B",X"0000",X"FFFA",X"FFFC",X"0002",X"0007",X"000A",X"FFFD",X"0006",X"FFFE",X"FFFD",X"0008",X"FFFD",X"FFFB",X"0003",X"FFF6",X"0000",X"FFFC",X"FFF5",X"0003",X"FFFA",X"FFFD",X"FFFF",X"FFF7",X"0005",X"FFFC",X"FFFC",X"000C",X"0000",X"000A",X"0000",X"0003",X"FFFE",X"FFFA",X"FFFC",X"000D",X"FFF8",X"FFFA",X"FFFE",X"0002",X"FFF5",X"0005",X"0005",X"FFF9",X"0000",X"0003",X"FFFA",X"FFFE",X"FFFD",X"0008",X"FFFC",X"FFF7",X"FFFE",X"0000",X"000D",X"FFF8",X"0007",X"FFFC",X"0003",X"FFFE",X"0001",X"0000",X"0003",X"FFFA",X"0000",X"0014",X"FFF7",X"0001",X"0000",X"0002",X"FFFF",X"0000",X"000B",X"0001",X"0008",X"0008",X"0000",X"FFFE",X"FFF8",X"0002",X"FFF4",X"0000",X"0000",X"FFF7",X"FFFD",X"FFFC",X"0000",X"FFF9",X"FFFF",X"FFFD",X"FFFC",X"0000",X"FFFE",X"FFFD",X"0007",X"0009",X"0000",X"FFF6",X"FFF8",X"FFF9",X"0000",X"0003",X"FFF8",X"FFFA",X"0000",X"FFF8",X"FFF6",X"FFFA",X"0007",X"0007",X"0008",X"000D",X"000F",X"000B",X"FFFE",X"0000",X"FFF4",X"0001",X"0000",X"0000",X"FFFD",X"000E",X"0004",X"0005",X"0002",X"000C",X"0007",X"FFF7",X"FFF8",X"FFF7",X"FFF7",X"FFFC",X"FFFF",X"FFFC",X"0002",X"0000",X"FFF0",X"0003",X"0008",X"0009",X"FFFC",X"0008",X"0007",X"0002",X"0006",X"FFFC",X"FFFB",X"FFF5",X"FFFB",X"0006",X"FFFD",X"FFF7",X"FFF7",X"0002",X"0003",X"FFFA",X"FFFB",X"FFFD",X"FFFF",X"0010",X"0005",X"0004",X"0004",X"FFFC",X"0006",X"FFFE",X"FFFB",X"0004",X"0001",X"000C",X"FFFF",X"FFFD",X"0008",X"FFFD",X"FFFE",X"0001",X"000A",X"0005",X"FFFF",X"FFF9",X"FFFB",X"0000",X"0000",X"0000",X"0001",X"0007",X"000C",X"FFFE",X"0007",X"FFFE",X"0000",X"0001",X"0002",X"FFFE",X"FFF6",X"0000",X"0008",X"FFF1",X"FFFF",X"0000",X"0001",X"FFFD",X"0000",X"0005",X"FFFC",X"0001",X"0000",X"FFFE",X"0000",X"0002",X"0000",X"0003",X"0002",X"0003",X"0000",X"FFFA",X"0005",X"0009",X"FFFA",X"FFFE",X"0005",X"0002",X"0006",X"FFFD",X"0006",X"FFFB",X"0000",X"0006",X"000A",X"FFFB",X"FFFD",X"0007",X"FFF9",X"FFFF",X"0003",X"0002",X"0002",X"FFFB",X"FFFA",X"0000",X"0000",X"FFFE",X"0007",X"0007",X"0001",X"FFFE",X"0009",X"0000",X"FFFF",X"0001",X"FFFD",X"FFF8",X"0001",X"0006",X"0000",X"0005",X"0005",X"0007",X"FFFB",X"FFF5",X"0000",X"FFFD",X"FFF5",X"FFF9",X"0008",X"0005",X"0000",X"0004",X"0006",X"FFFF",X"FFFC",X"FFFD",X"FFF8",X"FFFC",X"FFFF",X"0007",X"0013",X"FFFA",X"0000",X"0006",X"0001",X"0000",X"FFFF",X"0003",X"0000",X"FFFF",X"FFF6",X"FFF8",X"FFF5",X"FFF9",X"FFFB",X"FFFD",X"0002",X"0001",X"0000",X"0005",X"0006",X"0000",X"FFFE",X"0002",X"0000",X"FFF4",X"FFF9",X"0001",X"FFFC",X"FFFC",X"0001",X"FFFF",X"0008",X"FFFD",X"FFF3",X"FFF7",X"0002",X"0007",X"FFF8",X"0001",X"FFF8",X"0002",X"0005",X"000F",X"0006",X"0009",X"0009",X"FFFF",X"0000",X"FFFF",X"0010",X"FFFF",X"FFF9",X"FFF1",X"FFF3",X"FFEF",X"FFFD",X"FFFD",X"0001",X"FFFE",X"0001",X"0006",X"FFFE",X"FFFF",X"FFFB",X"0002",X"0000",X"0000",X"FFFE",X"FFF9",X"0001",X"0000",X"0010",X"0005",X"0001",X"FFFB",X"FFFC",X"0003",X"FFFC",X"FFF8",X"0002",X"0001",X"FFFF",X"0001",X"0006",X"0000",X"FFFB",X"FFFF",X"FFFB",X"FFF4",X"0008",X"FFFA",X"0003",X"0006",X"0001",X"FFF7",X"000A",X"FFFE",X"0002",X"FFFF",X"0008",X"0001",X"0003",X"0006",X"FFFF",X"0007",X"0000",X"0002",X"FFFD",X"FFFB",X"0002",X"FFFF",X"0000",X"FFFA",X"FFFC",X"000B",X"FFFA",X"FFF9",X"FFF4",X"FFF6",X"0006",X"0001",X"FFFF",X"FFFB",X"FFFC",X"0000",X"0000",X"0003",X"0005",X"0005",X"000F",X"FFFC",X"FFFB",X"FFFE",X"0000",X"0005",X"0007",X"0000",X"FFFD",X"0001",X"FFFC",X"FFF8",X"FFFE",X"FFFD",X"0009",X"FFFD",X"000B",X"0002",X"0002",X"FFFC",X"FFF6",X"FFF9",X"FFFD",X"FFFF",X"FFF5",X"FFFB",X"FFFD",X"FFFE",X"FFF8",X"FFFC",X"0000",X"FFFE",X"0000",X"0001",X"FFFD",X"FFFD",X"0002",X"0009",X"0007",X"0001",X"FFFD",X"0000",X"FFFD",X"0000",X"FFFE",X"0002",X"FFF7",X"FFFB",X"FFF1",X"FFFD",X"0000",X"FFFE",X"FFFC",X"FFF8",X"0001",X"0000",X"0005",X"FFFD",X"FFFA",X"0002",X"0007",X"FFF8",X"FFFE",X"0004",X"FFF7",X"0002",X"0009",X"FFFE",X"FFF4",X"FFFC",X"FFF9",X"FFF8",X"FFFA",X"0005",X"0009",X"FFFC",X"FFF6",X"FFFF",X"FFF4",X"FFFC",X"FFFD",X"0007",X"FFFD",X"0006",X"0000",X"FFFE",X"0006",X"0003",X"0000",X"0003",X"FFFD",X"FFFE",X"0001",X"FFFB",X"0000",X"0000",X"0004",X"FFF3",X"FFF9",X"FFFA",X"FFF3",X"0002",X"0005",X"0003",X"0009",X"FFFF",X"0000",X"FFF4",X"0000",X"0003",X"0008",X"0002",X"FFFC",X"0001",X"FFFF",X"0007",X"0002",X"0000",X"0013",X"FFF8",X"0009",X"0013",X"0008",X"0001",X"FFFA",X"0000",X"0000",X"FFFF",X"0000",X"0000",X"FFEB",X"0000",X"FFFD",X"0000",X"FFFA",X"0008",X"FFFA",X"0000",X"0004",X"0000",X"0009",X"0000",X"FFFB",X"FFFD",X"0000",X"FFFE",X"0000",X"0004",X"000A",X"0003",X"FFFF",X"FFFF",X"FFF6",X"FFFB",X"FFF6",X"0000",X"FFF8",X"0003",X"0002",X"0003",X"0007",X"FFFD",X"FFF8",X"0000",X"0001",X"FFFA",X"FFFC",X"FFFC",X"0000",X"0002",X"0008",X"FFFA",X"0006",X"000D",X"0009",X"0000",X"FFFF",X"FFF7",X"FFF4",X"0004",X"FFFA",X"FFF8",X"FFFC",X"0006",X"FFFF",X"FFF5",X"0001",X"0007",X"0001",X"FFF8",X"FFF8",X"0002",X"0001",X"0002",X"FFFE",X"0002",X"0002",X"0007",X"0000",X"0000",X"0008",X"0007",X"0000",X"FFFD",X"FFFA",X"FFFC",X"FFF9",X"0000",X"FFFD",X"000E",X"0003",X"FFFE",X"FFFD",X"0006",X"FFFE",X"0004",X"FFFB",X"0004",X"0006",X"0000",X"0003",X"0002",X"0001",X"0000",X"0002",X"0006",X"0005",X"0001",X"0000",X"0002",X"FFFE",X"FFFC",X"FFFB",X"0001",X"000B",X"0000",X"000B",X"0000",X"FFF4",X"FFFC",X"0000",X"FFFB",X"FFFD",X"000D",X"0009",X"0007",X"000D",X"0000",X"0009",X"0007",X"0000",X"FFF8",X"FFFB",X"FFF9",X"FFF4",X"FFF6",X"FFF8",X"0006",X"FFFF",X"FFFC",X"FFF6",X"000D",X"0005",X"0002",X"0001",X"0000",X"FFFD",X"0003",X"0001",X"0009",X"FFFC",X"0006",X"0007",X"0000",X"0003",X"FFFF",X"FFFC",X"FFF7",X"FFFD",X"0007",X"0000",X"0004",X"0004",X"FFF4",X"FFFA",X"0000",X"FFFF",X"0000",X"0000",X"0006",X"0000",X"0005",X"FFF4",X"0001",X"0003",X"000C",X"000C",X"0003",X"000A",X"0001",X"FFFD",X"0000",X"FFFE",X"FFF8",X"FFFD",X"0005",X"0001",X"FFF3",X"0004",X"0002",X"0004",X"0003",X"FFF8",X"FFF7",X"FFFB",X"0002",X"0008",X"0005",X"FFFA",X"0000",X"0004",X"0005",X"0000",X"FFFF",X"FFFC",X"FFFA",X"0000",X"FFFD",X"FFFE",X"0000",X"0001",X"000A",X"FFFC",X"0004",X"FFFE",X"FFF9",X"FFFB",X"0003",X"FFFF",X"0006",X"0008",X"0008",X"0000",X"0001",X"FFF9",X"0000",X"FFFF",X"FFF9",X"FFFB",X"FFFC",X"FFF0",X"0000",X"FFFE",X"0001",X"0008",X"FFFD",X"FFFE",X"0009",X"0003",X"FFFA",X"FFFE",X"FFFD",X"FFFC",X"0007",X"FFFD",X"0001",X"0005",X"0002",X"FFF5",X"FFFC",X"FFF8",X"FFF5",X"FFFD",X"0001",X"000C",X"000A",X"0001",X"0004",X"0000",X"FFFE",X"FFFD",X"0008",X"0003",X"0004",X"FFFA",X"FFEE",X"FFF4",X"0009",X"0005",X"0005",X"FFFF",X"FFF5",X"FFF6",X"0000",X"FFFD",X"FFF7",X"FFF7",X"0000",X"FFF9",X"FFF8",X"FFFB",X"FFF5",X"0000",X"FFFC",X"FFF9",X"FFFF",X"0008",X"0008",X"0005",X"0002",X"0003",X"0002",X"0009",X"FFFA",X"0004",X"FFFB",X"0004",X"0006",X"FFFD",X"0008",X"0008",X"FFFD",X"000A",X"FFFA",X"FFF8",X"FFFE",X"FFF9",X"FFF9",X"FFEC",X"FFF8",X"FFFA",X"0000",X"0001",X"FFFF",X"FFFB",X"0002",X"FFF6",X"0004",X"FFFF",X"0001",X"FFFB",X"0004",X"0010",X"0008",X"0004",X"0000",X"FFF7",X"0007",X"0000",X"FFFC",X"FFF1",X"FFF6",X"FFF9",X"FFFE",X"FFFC",X"000C",X"0001",X"0001",X"0000",X"FFFB",X"FFFB",X"0001",X"FFFE",X"FFFC",X"FFFD",X"0001",X"0000",X"FFF7",X"0001",X"0000",X"0007",X"0002",X"FFF5",X"0004",X"0005",X"0009",X"0000",X"0000",X"FFFD",X"FFFF",X"FFFD",X"0004",X"FFF1",X"FFF6",X"0000",X"FFF9",X"FFFF",X"FFF9",X"FFF5",X"0000",X"FFFE",X"FFFE",X"0006",X"0005",X"FFFC",X"FFF8",X"0004",X"FFFF",X"0002",X"0001",X"000A",X"0005",X"FFFC",X"0000",X"0003",X"0008",X"0000",X"FFF9",X"FFFF",X"0000",X"0002",X"FFF6",X"FFFE",X"0007",X"0005",X"FFFF",X"FFFD",X"0001",X"FFFD",X"FFF6",X"0001",X"0002",X"0003",X"0009",X"0001",X"FFF7",X"FFFC",X"0000",X"0000",X"0006",X"0004",X"0009",X"FFFA",X"0006",X"0003",X"FFFF",X"FFFF",X"FFFB",X"FFF8",X"FFF3",X"FFFA",X"FFFF",X"FFFF",X"0002",X"0007",X"0008",X"FFF8",X"FFFC",X"FFF7",X"0000",X"0005",X"0003",X"FFF6",X"0005",X"0008",X"000A",X"0007",X"0000",X"FFFF",X"0002",X"0004",X"FFF9",X"000A",X"FFF9",X"FFF6",X"FFED",X"FFF0",X"FFFD",X"FFF2",X"FFFF",X"0006",X"0007",X"FFFF",X"FFF8",X"FFFF",X"FFFD",X"FFFE",X"0004",X"0007",X"0005",X"0008",X"FFFA",X"0002",X"0005",X"FFFD",X"FFFF",X"0009",X"FFFB",X"FFF5",X"0004",X"0002",X"FFFF",X"FFF2",X"0001",X"0000",X"FFF5",X"FFFF",X"FFFC",X"FFF5",X"FFF5",X"FFF9",X"FFFC",X"000C",X"0008",X"0000",X"0004",X"FFFA",X"0001",X"0008",X"0000",X"FFFD",X"FFFC",X"FFFA",X"FFFB",X"FFFF",X"0006",X"0009",X"000A",X"0000",X"FFFF",X"FFFB",X"FFFD",X"FFFD",X"FFF2",X"FFF5",X"0000",X"0003",X"FFF2",X"FFFB",X"0000",X"0002",X"FFFF",X"FFFD",X"0003",X"0004",X"0000",X"0000",X"0000",X"0000",X"FFFA",X"FFFF",X"FFFF",X"000C",X"0001",X"0002",X"000C",X"FFF8",X"0000",X"0004",X"FFF9",X"FFFE",X"0008",X"FFFA",X"0000",X"0004",X"FFFB",X"FFFC",X"FFF9",X"FFFB",X"0001",X"FFFC",X"FFF0",X"0007",X"FFFD",X"000D",X"0001",X"FFFC",X"0005",X"FFFD",X"FFFE",X"FFFD",X"0003",X"0000",X"FFFD",X"0007",X"0003",X"FFF6",X"0000",X"0000",X"FFFF",X"0004",X"FFF9",X"FFFE",X"FFF7",X"FFF4",X"FFF6",X"FFF9",X"FFF7",X"FFF7",X"FFFC",X"0000",X"000B",X"FFFF",X"0001",X"0010",X"0007",X"0002",X"FFFC",X"0000",X"0008",X"FFFD",X"FFFE",X"FFF9",X"FFFF",X"FFF8",X"FFFB",X"FFFE",X"000A",X"0001",X"0000",X"FFFA",X"0000",X"FFFF",X"0001",X"FFFA",X"FFF8",X"0005",X"FFFD",X"FFF5",X"FFFD",X"0003",X"FFFB",X"0002",X"FFFB",X"0008",X"0003",X"FFFF",X"FFF5",X"FFFB",X"0003",X"0000",X"0000",X"0001",X"0000",X"FFFC",X"FFF8",X"0002",X"0001",X"0003",X"0003",X"0000",X"0009",X"FFFA",X"FFFC",X"FFF2",X"FFE9",X"FFF7",X"FFFC",X"FFF6",X"FFFE",X"0006",X"0008",X"000E",X"000C",X"FFFC",X"FFFF",X"FFFD",X"FFFC",X"0002",X"0012",X"0009",X"0009",X"0003",X"0005",X"FFF9",X"FFFE",X"FFEC",X"FFF0",X"FFF0",X"0000",X"0006",X"0000",X"FFF3",X"FFF9",X"FFFC",X"0004",X"0004",X"000C",X"000D",X"0009",X"0002",X"FFFD",X"FFF3",X"FFF7",X"0000",X"0001",X"0004",X"FFFA",X"0000",X"FFFD",X"FFFA",X"FFFF",X"0001",X"000B",X"0002",X"0006",X"0000",X"FFFE",X"0002",X"0003",X"FFFC",X"FFFF",X"FFFC",X"0004",X"FFFD",X"FFFA",X"0005",X"0002",X"0008",X"0000",X"FFFC",X"FFFB",X"FFF9",X"0009",X"FFFA",X"0004",X"FFF9",X"0000",X"0008",X"0000",X"0001",X"FFFC",X"0005",X"0001",X"0006",X"FFFC",X"0000",X"0000",X"0001",X"FFFA",X"000F",X"0005",X"000E",X"0001",X"0006",X"0005",X"FFFE",X"FFFC",X"FFFB",X"0007",X"FFFD",X"FFF5",X"FFF3",X"0001",X"FFFE",X"FFFD",X"0003",X"FFFE",X"0006",X"0000",X"0001",X"FFFC",X"FFF5",X"0003",X"FFFE",X"FFFC",X"FFFE",X"0000",X"0000",X"0000",X"0001",X"FFFF",X"FFFC",X"FFFF",X"FFFD",X"000B",X"0005",X"FFF5",X"FFF7",X"FFFB",X"FFFE",X"0000",X"FFFC",X"FFFD",X"0003",X"0004",X"FFFF",X"000E",X"FFF7",X"0004",X"0001",X"0009",X"0009",X"FFFE",X"0004",X"FFFB",X"FFF9",X"FFFC",X"FFF7",X"FFFD",X"0006",X"0000",X"FFF9",X"0001",X"FFF6",X"FFFB",X"FFF5",X"0000",X"0000",X"0001",X"0003",X"0008",X"000B",X"0009",X"FFF6",X"0006",X"FFFA",X"FFFE",X"FFF9",X"0007",X"FFFC",X"0005",X"0010",X"0004",X"0002",X"FFF8",X"FFFD",X"FFFE",X"FFF5",X"0000",X"0002",X"0002",X"FFFD",X"0003",X"FFFC",X"FFFE",X"000A",X"FFFE",X"FFF5",X"FFF8",X"FFF2",X"0004",X"0000",X"0009",X"FFFD",X"FFFA",X"0002",X"FFFB",X"0005",X"0000",X"FFFB",X"FFF6",X"0000",X"0004",X"FFFB",X"0000",X"0008",X"000B",X"0003",X"0006",X"FFFA",X"000A",X"FFFF",X"FFFF",X"0002",X"FFF5",X"FFFA",X"FFF5",X"FFFB",X"FFFD",X"FFFF",X"FFF8",X"FFFC",X"FFFA",X"FFFC",X"FFFF",X"0001",X"0004",X"0005",X"0003",X"0005",X"FFFD",X"0005",X"0005",X"FFFE",X"0003",X"0000",X"0000",X"FFFA",X"FFF9",X"FFFB",X"FFFB",X"FFFC",X"000D",X"FFFD",X"FFFF",X"FFF9",X"FFFF",X"FFFC",X"0000",X"0007",X"0003",X"0008",X"000C",X"0000",X"0008",X"0003",X"0002",X"0003",X"FFFC",X"0000",X"0006",X"0001",X"0003",X"0006",X"0009",X"0005",X"FFFB",X"0000",X"FFF9",X"FFF4",X"FFF9",X"0008",X"0004",X"0000",X"FFF6",X"0000",X"FFF6",X"0000",X"FFF8",X"FFF5",X"0001",X"0003",X"0007",X"FFFA",X"FFFE",X"FFFE",X"0002",X"0000",X"0007",X"0000",X"FFFF",X"0000",X"0004",X"FFFC",X"0000",X"FFFD",X"FFFD",X"FFFC",X"000F",X"FFF9",X"0000",X"0010",X"FFFD",X"0004",X"0009",X"FFFE",X"FFF8",X"0000",X"0001",X"FFFE",X"FFF7",X"FFF8",X"FFFF",X"0000",X"FFFA",X"FFF8",X"0000",X"0000",X"0006",X"FFF8",X"000B",X"000E",X"0007",X"0004",X"0001",X"0004",X"0004",X"000D",X"0003",X"0000",X"FFFE",X"0002",X"FFF4",X"0000",X"FFF8",X"FFFA",X"0001",X"0003",X"0003",X"0006",X"0008",X"FFFB",X"0003",X"0000",X"FFFA",X"FFFA",X"0005",X"000A",X"FFFB",X"FFFA",X"0003",X"0008",X"0005",X"0007",X"0007",X"FFFE",X"0002",X"FFFA",X"0005",X"0000",X"FFFF",X"0005",X"FFF9",X"FFFF",X"0000",X"0008",X"0009",X"0001",X"FFFB",X"0002",X"FFF6",X"0008",X"FFF8",X"FFFE",X"FFF1",X"0000",X"0000",X"FFFD",X"FFF4",X"FFF7",X"0003",X"0001",X"0000",X"0007",X"0008",X"0003",X"0006",X"FFFD",X"FFFF",X"FFFA",X"0007",X"0004",X"0007",X"000D",X"000C",X"FFF9",X"FFF4",X"FFF7",X"FFF9",X"0008",X"FFF3",X"FFFE",X"0000",X"FFF2",X"0000",X"0004",X"FFFC",X"000E",X"0001",X"0005",X"FFFE",X"FFF8",X"FFFD",X"0000",X"FFFD",X"FFFA",X"FFFE",X"0000",X"0002",X"0006",X"000B",X"FFFF",X"0003",X"0002",X"FFFE",X"FFFD",X"0005",X"0006",X"0005",X"0002",X"FFFD",X"FFFC",X"FFFB",X"0000",X"0006",X"0000",X"0002",X"FFFE",X"FFFB",X"FFFD",X"FFF6",X"FFF3",X"FFF9",X"FFFB",X"0001",X"0003",X"FFFF",X"FFFB",X"0013",X"000D",X"FFFE",X"0000",X"0001",X"FFFB",X"FFFB",X"FFFC",X"0000",X"FFFD",X"0004",X"0001",X"FFFE",X"0001",X"0005",X"FFF9",X"0003",X"0001",X"FFF8",X"FFF4",X"FFFD",X"FFF7",X"0009",X"0006",X"0004",X"0009",X"000B",X"0004",X"0000",X"0003",X"0000",X"0002",X"0004",X"FFF6",X"FFF8",X"FFEC",X"FFFA",X"0004",X"0001",X"0007",X"FFF9",X"FFFC",X"0000",X"FFFE",X"FFFB",X"FFFD",X"0001",X"000D",X"000C",X"0008",X"000B",X"0001",X"0000",X"FFFD",X"FFFC",X"FFFD",X"0004",X"0002",X"FFFC",X"0000",X"FFFD",X"FFFE",X"0000",X"FFFA",X"FFFC",X"FFF5",X"FFFA",X"0008",X"0005",X"0002",X"0003",X"FFF4",X"FFFB",X"0003",X"FFFF",X"FFFC",X"0005",X"FFFB",X"0004",X"0000",X"FFFE",X"0007",X"FFFB",X"0002",X"0005",X"0001",X"FFFB",X"0005",X"0000",X"FFFD",X"FFFD",X"FFFE",X"FFF8",X"FFF9",X"0003",X"0001",X"0000",X"0002",X"0012",X"FFFC",X"FFF7",X"0000",X"FFFB",X"FFFF",X"FFFA",X"0001",X"FFF9",X"FFFC",X"FFFC",X"FFFE",X"FFFE",X"FFFA",X"0000",X"FFFA",X"FFFA",X"0009",X"0001",X"FFFD",X"0002",X"0002",X"FFF9",X"FFF3",X"0003",X"0006",X"0002",X"0007",X"0004",X"FFFF",X"0004",X"0005",X"0003",X"0000",X"000A",X"0006",X"FFF6",X"0001",X"FFF6",X"0007",X"FFFB",X"0002",X"FFFB",X"FFF9",X"FFF7",X"FFFA",X"FFFF",X"0009",X"0005",X"0009",X"0006",X"0009",X"0003",X"0000",X"FFFF",X"0000",X"FFFC",X"FFFE",X"FFFB",X"0001",X"FFFC",X"FFF9",X"FFFD",X"FFF8",X"FFFD",X"0000",X"FFFC",X"FFFC",X"0003",X"0004",X"0009",X"0002",X"0006",X"FFF7",X"FFFB",X"0003",X"FFFC",X"0001",X"FFF2",X"FFFA",X"000A",X"0000",X"0001",X"0008",X"0001",X"FFF7",X"0001",X"0002",X"FFF8",X"FFF7",X"FFFC",X"000E",X"0005",X"0002",X"FFFD",X"FFFC",X"FFFC",X"0002",X"FFF5",X"FFF8",X"0001",X"0004",X"0000",X"0010",X"FFFA",X"0000",X"FFFA",X"FFFD",X"FFFD",X"FFF8",X"0003",X"FFFB",X"000C",X"0012",X"0000",X"FFFA",X"FFFD",X"FFFC",X"FFFF",X"FFFF",X"FFFC",X"FFFE",X"FFFA",X"FFFD",X"FFFF",X"FFFF",X"0001",X"0001",X"FFFB",X"0000",X"0005",X"FFFC",X"FFF8",X"FFF9",X"FFFE",X"0005",X"0003",X"0006",X"000A",X"0005",X"0006",X"000A",X"FFFB",X"FFFF",X"0007",X"0000",X"0000",X"0000",X"FFF6",X"FFF9",X"FFF9",X"FFFD",X"0005",X"0005",X"0000",X"FFF5",X"FFF5",X"FFF6",X"FFFD",X"0007",X"000C",X"0008",X"0003",X"0014",X"0005",X"0002",X"FFFE",X"FFF6",X"0004",X"0004",X"0007",X"FFFD",X"FFFF",X"FFFB",X"0001",X"0004",X"FFF9",X"FFF7",X"FFFE",X"FFF3",X"FFFC",X"FFF5",X"0000",X"FFFD",X"0009",X"0000",X"000D",X"FFFE",X"0000",X"0000",X"0000",X"0000",X"FFFD",X"FFFB",X"0001",X"0006",X"0009",X"0002",X"FFFE",X"0003",X"FFF4",X"FFFD",X"000E",X"FFFE",X"0000",X"0008",X"0001",X"000B",X"0000",X"0004",X"FFFB",X"FFFF",X"000A",X"FFFE",X"FFF7",X"FFFD",X"FFF8",X"0006",X"0002",X"0000",X"0003",X"0000",X"FFFC",X"FFFC",X"FFFC",X"FFFB",X"0000",X"0008",X"000B",X"FFF9",X"0002",X"0006",X"0001",X"FFFB",X"FFF7",X"FFF6",X"FFF4",X"FFFB",X"FFFC",X"000D",X"0006",X"0001",X"0004",X"FFF9",X"0000",X"0000",X"0002",X"0003",X"FFFE",X"FFF8",X"0008",X"FFFA",X"0002",X"FFFC",X"FFFA",X"0005",X"0004",X"FFFA",X"FFFA",X"FFEC",X"FFF3",X"FFF4",X"FFF1",X"FFFE",X"000B",X"0004",X"0008",X"000B",X"0004",X"0006",X"0000",X"0009",X"0006",X"FFF9",X"FFFC",X"0004",X"FFFF",X"FFFB",X"0002",X"FFFC",X"FFFD",X"0001",X"0000",X"0005",X"0001",X"FFFB",X"0001",X"FFFC",X"FFFC",X"FFFC",X"0008",X"0000",X"FFFB",X"0003",X"0008",X"0004",X"0005",X"0004",X"FFF9",X"FFF5",X"FFFF",X"0002",X"FFF9",X"FFFB",X"0002",X"0003",X"0005",X"0000",X"FFF9",X"0004",X"0004",X"FFF8",X"FFF0",X"FFF9",X"FFF7",X"FFF3",X"FFF8",X"0009",X"000C",X"FFFD",X"0001",X"0003",X"0000",X"000C",X"0005",X"0004",X"0005",X"FFFE",X"FFFE",X"0008",X"0001",X"FFF9",X"0008",X"0004",X"0005",X"FFF7",X"FFF5",X"FFEF",X"FFF6",X"FFFA",X"FFFA",X"0006",X"0003",X"FFFC",X"0005",X"FFFE",X"FFFD",X"0000",X"0000",X"FFF2",X"FFFE",X"0000",X"FFFF",X"0000",X"FFFB",X"FFFC",X"0006",X"0001",X"FFFF",X"000D",X"000A",X"FFF8",X"0001",X"FFFC",X"0008",X"FFF8",X"0006",X"FFFF",X"0000",X"0007",X"FFFF",X"FFF7",X"0007",X"0006",X"FFF4",X"FFF4",X"FFF8",X"FFFB",X"0000",X"FFF8",X"FFF7",X"FFF9",X"FFFE",X"FFFF",X"FFFF",X"0000",X"0004",X"FFFB",X"0008",X"FFFF",X"0004",X"FFFC",X"FFFD",X"0000",X"0008",X"0004",X"000A",X"0007",X"000F",X"0001",X"FFF5",X"0002",X"0002",X"FFFB",X"0000",X"0000",X"0005",X"0001",X"FFF4",X"0000",X"FFF4",X"FFF2",X"FFFD",X"FFF9",X"FFF7",X"0004",X"0005",X"0002",X"0004",X"FFFE",X"0006",X"0000",X"0007",X"0009",X"0001",X"0002",X"0005",X"0008",X"FFFE",X"FFF8",X"FFF7",X"0000",X"FFF7",X"FFFA",X"0004",X"0003",X"0001",X"FFFE",X"0006",X"FFFC",X"0002",X"000D",X"FFFC",X"0002",X"FFF9",X"0000",X"0000",X"FFFF",X"0005",X"0001",X"FFFF",X"FFF8",X"0000",X"FFFF",X"FFEE",X"FFF6",X"FFF2",X"0002",X"FFFF",X"FFFD",X"FFFB",X"0001",X"0008",X"0006",X"0005",X"0004",X"0000",X"FFF5",X"0007",X"0009",X"FFFB",X"0000",X"0008",X"0000",X"FFF9",X"0000",X"FFF7",X"0000",X"0000",X"FFFE",X"0000",X"FFF7",X"FFF8",X"FFFC",X"0001",X"FFFE",X"FFF6",X"FFFB",X"FFFB",X"FFFA",X"FFF8",X"FFF0",X"FFFC",X"0000",X"000B",X"000F",X"0004",X"0000",X"0001",X"FFFC",X"000E",X"FFF7",X"FFF9",X"0005",X"FFFB",X"0003",X"0001",X"FFF8",X"FFF8",X"FFF7",X"FFF9",X"FFF9",X"FFFA",X"0001",X"0000",X"0003",X"0000",X"FFFF",X"0000",X"0004",X"FFF8",X"0008",X"0005",X"FFF8",X"0004",X"FFFC",X"0004",X"FFFA",X"FFFA",X"0001",X"FFFE",X"0007",X"0000",X"0003",X"0000",X"0001",X"FFFE",X"FFF7",X"FFF0",X"0000",X"0007",X"0002",X"FFFB",X"0000",X"0008",X"0002",X"FFFC",X"FFFE",X"FFFD",X"0002",X"0003",X"0002",X"FFFB",X"0003",X"0001",X"0003",X"0000",X"000B",X"FFF8",X"FFF5",X"0004",X"000B",X"0006",X"0003",X"FFFB",X"FFF1",X"FFFF",X"0010",X"FFFE",X"0005",X"FFF8",X"FFF6",X"FFFE",X"0000",X"0008",X"FFFB",X"0004",X"0000",X"0001",X"FFFF",X"FFFA",X"0000",X"FFF5",X"FFFB",X"0001",X"FFF8",X"FFFD",X"FFFC",X"000F",X"FFFF",X"FFFF",X"0000",X"FFFD",X"0002",X"0000",X"0004",X"0000",X"FFFA",X"FFFD",X"FFFA",X"000B",X"0008",X"0007",X"000E",X"0000",X"FFF6",X"0000",X"0007",X"FFFE",X"0004",X"FFFB",X"FFFE",X"FFF7",X"FFF9",X"FFFE",X"0006",X"0007",X"FFFF",X"0000",X"FFF6",X"0000",X"FFFD",X"0003",X"0001",X"0008",X"0003",X"FFF9",X"000A",X"0009",X"000B",X"0007",X"0008",X"0003",X"FFF8",X"FFF8",X"FFF5",X"FFFE",X"0008",X"FFF6",X"0001",X"0001",X"FFF9",X"FFFB",X"FFFD",X"0000",X"0003",X"0000",X"0000",X"0002",X"0001",X"FFFF",X"0009",X"0005",X"FFFC",X"FFF9",X"FFF3",X"0001",X"FFFF",X"FFF6",X"FFED",X"FFF5",X"FFFD",X"0003",X"000E",X"FFFA",X"0007",X"FFFA",X"0000",X"0009",X"0000",X"0000",X"FFF3",X"FFFA",X"FFF1",X"0002",X"FFF6",X"FFFD",X"FFFE",X"FFFA",X"0002",X"0003",X"0005",X"FFFD",X"FFFE",X"FFFF",X"0000",X"0001",X"FFFB",X"FFFD",X"0001",X"0001",X"0004",X"FFF8",X"0000",X"0014",X"000B",X"000C",X"FFF9",X"FFFE",X"0004",X"FFFF",X"0000",X"0006",X"0005",X"0000",X"FFFA",X"FFFB",X"000C",X"0001",X"FFFD",X"0000",X"0006",X"000A",X"FFFF",X"FFFD",X"0004",X"0001",X"0008",X"0000",X"FFFB",X"FFF3",X"FFFF",X"FFF4",X"FFEF",X"0006",X"0000",X"0005",X"0006",X"FFFF",X"FFFE",X"0001",X"000B",X"0005",X"FFFF",X"0000",X"FFFE",X"FFF7",X"FFF8",X"FFFD",X"0003",X"0005",X"0005",X"0000",X"FFF7",X"FFF6",X"FFF4",X"0006",X"0000",X"0002",X"0003",X"FFFE",X"FFFD",X"FFF6",X"0001",X"0006",X"0004",X"FFFE",X"0000",X"FFFE",X"0004",X"0007",X"0001",X"FFFC",X"FFFF",X"0002",X"0004",X"FFF9",X"0005",X"0005",X"0000",X"0001",X"FFFD",X"FFFE",X"0000",X"0001",X"FFF6",X"FFFC",X"0007",X"FFFE",X"0000",X"000A",X"0002",X"0002",X"0000",X"0001",X"FFF8",X"FFFD",X"0007",X"FFF2",X"FFF7",X"FFF7",X"FFFB",X"FFFA",X"0001",X"0000",X"0002",X"0009",X"FFFC",X"0004",X"0007",X"0004",X"0009",X"FFFA",X"0003",X"FFF8",X"0001",X"0003",X"0004",X"0008",X"0000",X"000C",X"0004",X"FFFE",X"FFF9",X"FFFB",X"0000",X"0001",X"FFFC",X"0001",X"FFF9",X"FFF7",X"0004",X"0001",X"0000",X"0009",X"FFFD",X"FFF5",X"FFF9",X"FFF8",X"0002",X"0000",X"FFFE",X"000C",X"000A",X"0003",X"FFFE",X"FFFC",X"0000",X"0004",X"0003",X"0000",X"0002",X"FFFE",X"FFF2",X"FFFF",X"000B",X"0007",X"FFFE",X"FFFE",X"FFFF",X"0007",X"0004",X"0007",X"0001",X"FFF3",X"FFEF",X"FFFC",X"FFFB",X"FFFE",X"FFF5",X"0004",X"FFF3",X"0001",X"0007",X"0002",X"0008",X"000C",X"000C",X"0008",X"0009",X"000C",X"0002",X"FFF8",X"0000",X"0001",X"FFF8",X"FFF9",X"FFF1",X"FFF8",X"FFF8",X"FFFD",X"FFFC",X"0003",X"FFFD",X"FFF9",X"0005",X"0000",X"FFF4",X"FFF5",X"0003",X"000F",X"0007",X"000C",X"0005",X"0001",X"0006",X"FFFB",X"FFF9",X"0000",X"FFFB",X"0000",X"0003",X"000A",X"0000",X"FFF9",X"0001",X"0002",X"FFFC",X"FFFD",X"0001",X"0009",X"FFF4",X"FFEF",X"FFF7",X"0009",X"0006",X"0017",X"0001",X"FFFE",X"0007",X"FFFE",X"000C",X"0005",X"0003",X"0003",X"FFFA",X"FFF5",X"FFF1",X"000B",X"0001",X"FFF5",X"000D",X"0001",X"0008",X"FFFD",X"0006",X"FFF8",X"FFF0",X"FFED",X"FFFB",X"FFF2",X"0000",X"0002",X"0005",X"0009",X"0003",X"FFFC",X"0006",X"0007",X"FFFD",X"0009",X"000B",X"0007",X"FFF2",X"FFFE",X"FFF7",X"FFFB",X"FFFE",X"FFF9",X"FFFA",X"0009",X"FFFE",X"FFF4",X"0005",X"0007",X"0000",X"FFFE",X"000B",X"0009",X"FFF9",X"FFF4",X"0003",X"FFF3",X"FFEA",X"FFF4",X"FFFE",X"0007",X"0007",X"0012",X"000E",X"0003",X"FFF8",X"0010",X"000A",X"FFF8",X"FFFB",X"0008",X"FFF9",X"FFED",X"FFF9",X"FFF2",X"0009",X"FFFB",X"000C",X"0019",X"0004",X"0002",X"0000",X"FFF8",X"0000",X"0009",X"FFF9",X"0005",X"0010",X"0000",X"0003",X"0004",X"0006",X"FFEE",X"FFFD",X"0004",X"FFF6",X"FFF1",X"0002",X"0005",X"0000",X"FFF3",X"0004",X"0015",X"0005",X"0002",X"000B",X"0007",X"0000",X"FFFC",X"0004",X"0003",X"FFF0",X"FFFB",X"0004",X"FFF5",X"FFFB",X"FFFC",X"0005",X"0000",X"000E",X"0018",X"000C",X"000C",X"FFF6",X"FFFA",X"FFFD",X"FFF6",X"FFFE",X"0008",X"0002",X"FFFF",X"FFFD",X"FFFE",X"0003",X"FFFE",X"0004",X"0011",X"0011",X"0003",X"FFFD",X"FFFC",X"FFF8",X"FFF6",X"0001",X"000B",X"FFE8",X"FFF2",X"FFFD",X"FFE1",X"FFDB",X"FFEB",X"FFF4",X"FFE6",X"FFEE",X"0006",X"0002",X"FFFD",X"002B",X"0029",X"002C",X"003F",X"0041",X"004A",X"003A",X"0057",X"004A",X"004F",X"0036",X"FEFD",X"FEA2",X"FFB9",X"FFFC",X"0024",X"FF92",X"FEC2",X"0166",X"0395",X"0310",X"0312",X"010D",X"00E1",X"FE2D",X"FA0C",X"F3E5",X"F06A",X"F607",X"F896",X"00B6",X"0E2F",X"1832",X"1B6E",X"1848",X"0F7A",X"FB61",X"EC13",X"E59D",X"E7EE",X"F1A2",X"F7CC",X"FCB5",X"0231",X"0B70",X"0DD0",X"0A94",X"0CDD",X"0BC6",X"0370",X"023C",X"02E3",X"FAF3",X"F0C3",X"E59D",X"E361",X"EFA3",X"F7FE",X"FFA3",X"09DA",X"18B1",X"1FED",X"1A52",X"1AD4",X"1A28",X"0889",X"F2F5",X"EE3C",X"ECE0",X"EA51",X"E211",X"D6C0",X"E186",X"F48A",X"067B",X"16E1",X"253B",X"2B34",X"2025",X"0FBA",X"052A",X"FE05",X"F178",X"EB63",X"F14F",X"F8A7",X"FA73",X"EAB5",X"E00E",X"E5A6",X"F215",X"01D5",X"174D",X"2B1C",X"2FDB",X"27EA",X"1C1B",X"0D82",X"F6CE",X"E1DA",X"E040",X"E661",X"EDDE",X"E68F",X"DA87",X"E6E7",X"FD87",X"0C5C",X"19E6",X"2C54",X"35C1",X"2A3D",X"146A",X"FE54",X"ED1F",X"DBE2",X"D82E",X"E704",X"FC88",X"031C",X"F06F",X"E918",X"F853",X"0476",X"073D",X"0F47",X"1E0A",X"22C0",X"1C30",X"0E90",X"008D",X"F491",X"EE53",X"F3B1",X"FCA1",X"0077",X"EEEE",X"DCB6",X"E7D9",X"FD25",X"02F9",X"040F",X"0F03",X"18DE",X"19CA",X"14BF",X"0C75",X"03F3",X"F841",X"F4D0",X"F8C0",X"FF3B",X"F661",X"DDC5",X"D878",X"EEB3",X"0287",X"066A",X"0D8C",X"1AC6",X"1F84",X"1BAE",X"1302",X"0B20",X"FF5F",X"F6FC",X"F3CE",X"F6A1",X"F98D",X"E85B",X"D5C5",X"E21A",X"FE13",X"09DB",X"0AEA",X"1346",X"17F0",X"170C",X"11FC",X"0A48",X"FF95",X"F7AC",X"F85B",X"FD41",X"072F",X"01E0",X"E7AD",X"DD04",X"EE38",X"FCB5",X"FB03",X"FFFE",X"0BA3",X"12D3",X"1597",X"13B0",X"0C4C",X"0067",X"FB30",X"FAB9",X"033E",X"0C04",X"FD18",X"E400",X"E3B1",X"F54A",X"F9AE",X"F875",X"0100",X"09AB",X"1068",X"139D",X"1434",X"0CFD",X"04B2",X"FDD0",X"FC2B",X"0835",X"0881",X"EDDF",X"D937",X"E1A5",X"EE10",X"F048",X"FBEA",X"0BDF",X"1832",X"1D0D",X"1E1B",X"1963",X"0D71",X"0003",X"F1C5",X"F43E",X"0315",X"FC17",X"E5B2",X"E42A",X"F584",X"F956",X"F86C",X"FEEA",X"07AD",X"0E8A",X"11B4",X"135B",X"0DBB",X"0719",X"FDF0",X"F9A6",X"0922",X"1153",X"FBF4",X"E4DE",X"E79D",X"ED9A",X"EB35",X"F0C4",X"FD39",X"0B13",X"126F",X"17AB",X"1578",X"0EC6",X"066E",X"F9E5",X"FDE0",X"1058",X"0C88",X"F138",X"E4A0",X"EBDB",X"EC8F",X"ECEF",X"F3F1",X"01A7",X"0D75",X"15D0",X"192E",X"14B9",X"0ED3",X"0277",X"F995",X"069D",X"1196",X"FE2C",X"E245",X"DFD3",X"E4C0",X"E574",X"EADF",X"F912",X"0AF7",X"187F",X"224A",X"219D",X"1AFE",X"0F2E",X"FC92",X"FA23",X"0A06",X"09A8",X"EED9",X"DEDB",X"E2E3",X"E5D8",X"E7FE",X"EF28",X"FEDE",X"0C70",X"1803",X"1D6B",X"19DF",X"1459",X"0631",X"F99A",X"0390",X"1213",X"0536",X"EB7F",X"E5F1",X"E89E",X"EA53",X"EC9E",X"F5F3",X"01A6",X"0C62",X"1675",X"1730",X"1477",X"0D47",X"FD31",X"FAB4",X"0D08",X"1287",X"F9CE",X"E6A4",X"E3F6",X"E5B7",X"E7CE",X"EF73",X"FDA6",X"0A3E",X"1700",X"1D2E",X"1C05",X"19B1",X"0BCE",X"FB22",X"FFBB",X"0F1A",X"0439",X"EA35",X"DECB",X"DD80",X"DEF9",X"E389",X"F110",X"01C0",X"1325",X"2282",X"2578",X"239C",X"1AE3",X"05D6",X"F984",X"04D0",X"098A",X"F2FD",X"DF37",X"DAC9",X"DF08",X"E51A",X"F137",X"01BC",X"108E",X"1ED5",X"2323",X"1EC8",X"193E",X"089C",X"F2DF",X"F281",X"0461",X"00C9",X"EE01",X"E40C",X"E665",X"EBE4",X"F227",X"FCEF",X"078A",X"130F",X"1C03",X"1ACC",X"17C5",X"1010",X"FBAC",X"ECC4",X"FAA7",X"082F",X"FD98",X"ED62",X"E7A3",X"EA9E",X"EE52",X"F510",X"FE4B",X"08DE",X"15F2",X"1B29",X"193D",X"16EE",X"0A42",X"F32A",X"F0C3",X"0468",X"0803",X"F9A1",X"ED81",X"EC1A",X"ED86",X"EF6A",X"F500",X"FB8F",X"06CC",X"1226",X"14F2",X"16E9",X"156A",X"048F",X"F370",X"FE89",X"0D27",X"072F",X"F70A",X"EE39",X"EC89",X"EADC",X"ED50",X"F29A",X"FB9F",X"0A8A",X"13D3",X"1739",X"1A8E",X"1468",X"FD8C",X"F6B5",X"054C",X"0A1E",X"FCBC",X"EE3F",X"EA74",X"EA32",X"EC48",X"F207",X"F8CC",X"0554",X"11E7",X"1692",X"18A4",X"1A7B",X"0A59",X"F5E2",X"FB38",X"085C",X"049F",X"F426",X"EA1F",X"E8BD",X"E9CD",X"EF96",X"F5DC",X"FE50",X"0BFA",X"1537",X"17E2",X"1C5E",X"1810",X"00E2",X"F5C2",X"00E7",X"0826",X"FD95",X"EEA9",X"E98F",X"E97F",X"EC60",X"F158",X"F5D5",X"00E4",X"0DC1",X"142E",X"18CB",X"1EDC",X"1107",X"FAA7",X"FA6F",X"0770",X"0802",X"F92F",X"ED4B",X"E940",X"E827",X"EBA8",X"EF3D",X"F7B8",X"068B",X"12B1",X"1739",X"1F3D",X"1E8E",X"0772",X"F719",X"FDDA",X"07CD",X"0092",X"F166",X"E977",X"E71C",X"EA3C",X"EF46",X"F470",X"FFB4",X"0E4A",X"14CC",X"1933",X"2143",X"158E",X"FDB6",X"F74C",X"0297",X"066B",X"F9D4",X"ED84",X"E8B4",X"E912",X"ED34",X"EFC7",X"F5EC",X"03A6",X"100B",X"14BA",X"1EB7",X"212B",X"0D7B",X"FA68",X"FC93",X"06C8",X"036C",X"F5FC",X"ECE0",X"E899",X"E9EB",X"EBD4",X"EE90",X"F810",X"07EE",X"100D",X"1727",X"2202",X"1AA7",X"03AF",X"F8A8",X"019E",X"0863",X"FF58",X"F375",X"EC01",X"EB2C",X"EDC5",X"EFB5",X"F2BF",X"FE78",X"0A22",X"0E79",X"1973",X"1FC9",X"10F2",X"FCA2",X"FAFB",X"062E",X"066B",X"FB70",X"F106",X"EBF9");

 
 begin

    if (resetN='0') then
		Q_tmp <= ( others => '0');
    elsif(rising_edge(CLK)) then
--      if (ENA='1') then
		Q_tmp <= sin_table(conv_integer(ADDR));
--      end if;
   end if;
  end process;
 Q <= Q_tmp; 

		   
end arch;