library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.std_logic_signed.all;
use ieee.numeric_std.all;
-- Alex Grinshpun July 24 2017 
-- Dudy Nov 13 2017


entity back_gr_note is
port 	(
	   CLK      : in std_logic;
		RESETn	: in std_logic;
		oCoord_X : in integer;
		oCoord_Y : in integer;
		make    : in std_logic_vector(12 downto 0);
		drawing_request	: out std_logic;
		mVGA_RGB	: out std_logic_vector(7 downto 0)
	);
end back_gr_note;

architecture arc_back_gr_note of back_gr_note is 

-- Constants for frame drawing
constant	x_frame	: integer :=	639;
constant	y_frame	: integer :=	479;
constant	pianoHight : integer := 100;
constant	note_width : integer := 46;

signal mVGA_R	: std_logic_vector(2 downto 0); --	,	 			//	VGA Red[2:0]
signal mVGA_G	: std_logic_vector(2 downto 0); --	,	 			//	VGA Green[2:0]
signal mVGA_B	: std_logic_vector(1 downto 0); --	,  			//	VGA Blue[1:0]

	
begin

mVGA_RGB <=  mVGA_R & mVGA_G &  mVGA_B ;
-- defining three rectangles 

process ( oCoord_X,oCoord_y )
begin 
	if oCoord_Y > y_frame - pianoHight then
		mVGA_R <= "000";
		mVGA_G <= "000";
		mVGA_B <= "00";
		for i in 0 to 4 loop
			if oCoord_X >=note_width*i +3*i and oCoord_X <= note_width*(i+1) +3*i then
				if make(i) = '1' then
						mVGA_R <= "111";
						mVGA_G <= "100";
						mVGA_B <= "00";
				elsif i = 0 or i = 2 or i = 4 then
						mVGA_R <= "111";
						mVGA_G <= "111";
						mVGA_B <= "11";
				end if;
			end if;
		end loop;
		for i in 5 to 11 loop
			if oCoord_X >=note_width*i + 3*i and oCoord_X <= note_width*(i+1) +3*i  then
				if make(i) = '1' then
					mVGA_R <= "111";
					mVGA_G <= "100";
					mVGA_B <= "00";
				elsif i = 5 or i = 7 or i = 9 or i = 11 then
						mVGA_R <= "111";
						mVGA_G <= "111";
						mVGA_B <= "11";
				end if;
			end if;
		end loop;
		if oCoord_X >=note_width*12 +36  and oCoord_X <= x_frame -3  then
			if make(12) = '1' then
				mVGA_R <= "111";
				mVGA_G <= "100";
				mVGA_B <= "00";
			else
				mVGA_R <= "111";
				mVGA_G <= "111";
				mVGA_B <= "11";
			end if;
		end if;
		drawing_request <= '1';
	else
		drawing_request <= '0';
	end if;
end process ; 	
end architecture;		