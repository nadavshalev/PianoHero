library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_signed.all ;
use ieee.std_logic_arith.all;
library work;
use work.pkg2.all;

entity wisle_effect is
port(
  CLK     					: in std_logic;
  resetN 					: in std_logic;
  addrArr    				: in Arr_type;
  Q       					: out std_logic_vector(15 downto 0)
);
end wisle_effect;

architecture arch of wisle_effect is
	constant array_size 			: integer := 3001 ;
	
	signal Q_tmp       			:  std_logic_vector(15 downto 0) ;
	
	type table_type is array(0 to array_size - 1) of std_logic_vector(15 downto 0);
	constant sound0 : table_type := (X"FFEF",X"FFCD",X"FFD4",X"FFF0",X"FFF0",X"FFF7",X"0000",X"002E",X"003F",X"0029",X"0025",X"FFE7",X"FFC8",X"FFD5",X"FFD7",X"FFA0",X"FF9D",X"FFA3",X"FF7D",X"FF86",X"FF8B",X"FF7C",X"FF75",X"FF66",X"FF75",X"FF98",X"FFBE",X"FFF8",X"000C",X"0037",X"FFF8",X"FFC7",X"FFC0",X"FFE0",X"000F",X"FFE3",X"FFDE",X"FFD8",X"FFE5",X"FFFF",X"FFDC",X"FFB3",X"FFCD",X"FFD6",X"FFB9",X"FFB6",X"FFB6",X"FFCD",X"FFB4",X"FFBA",X"FFC6",X"FFED",X"000D",X"0017",X"0026",X"0040",X"0054",X"004C",X"0054",X"0022",X"000E",X"0015",X"0013",X"FFDD",X"FFC6",X"FFDA",X"FFE5",X"FFBF",X"FFB8",X"FFE0",X"FFE0",X"0006",X"FFFF",X"0001",X"0018",X"0044",X"0074",X"0096",X"0055",X"005B",X"0046",X"006E",X"0068",X"003F",X"0037",X"002E",X"002E",X"002E",X"0027",X"0024",X"0023",X"0047",X"005F",X"007D",X"0082",X"0080",X"007E",X"0096",X"0098",X"0077",X"009C",X"00CB",X"00C4",X"00AF",X"0095",X"0083",X"0062",X"002D",X"0028",X"003A",X"0017",X"FFFF",X"FFDB",X"FFB2",X"FFC2",X"FFDA",X"FFE2",X"FFE4",X"FFC7",X"FFDD",X"FFF5",X"FFED",X"FFCF",X"FFBA",X"FFC6",X"0006",X"0027",X"0029",X"0022",X"0020",X"0040",X"003E",X"0056",X"005C",X"0057",X"004F",X"0022",X"FFFF",X"FFE7",X"FF68",X"FF20",X"FF28",X"FEE1",X"FEF5",X"FEFE",X"FF08",X"FF35",X"FF6C",X"FFA8",X"FF7E",X"FF69",X"FF8C",X"FF9D",X"FF88",X"FF7A",X"FF82",X"FF57",X"FF3D",X"FF1F",X"FF06",X"FEFE",X"FF40",X"FF90",X"FFB2",X"FF90",X"FF73",X"FF9F",X"FFD0",X"FFE5",X"FFE6",X"FFFA",X"0018",X"004C",X"009F",X"0084",X"006E",X"0062",X"0042",X"0043",X"FFED",X"FFC4",X"FFD4",X"FFEE",X"FFFB",X"FFFE",X"FFDE",X"FFEA",X"FFEE",X"FFE7",X"FFCE",X"FFF6",X"FFFE",X"0007",X"001C",X"0037",X"0007",X"FFFD",X"000B",X"0076",X"00BD",X"00F2",X"0101",X"00EC",X"0092",X"0035",X"002E",X"000C",X"FFC3",X"FFA6",X"FF5B",X"FF3A",X"FF17",X"FF24",X"FF05",X"FECF",X"FEED",X"FF57",X"FFA6",X"FFD8",X"FFDF",X"FF9F",X"FFAD",X"FFA5",X"FFFD",X"002D",X"0072",X"0044",X"0020",X"0000",X"FFF4",X"FFD9",X"0031",X"0061",X"0057",X"003D",X"009F",X"0095",X"00BC",X"00E7",X"00E5",X"00CF",X"00B1",X"0086",X"0072",X"0034",X"0013",X"FFFB",X"FFDB",X"FFBE",X"FFF9",X"FFFA",X"FFF1",X"FFEF",X"FFED",X"000A",X"0044",X"0005",X"FFE4",X"FFFD",X"FFF9",X"FFED",X"FFEA",X"0031",X"0040",X"007A",X"00A1",X"00CC",X"00D7",X"0147",X"0191",X"0193",X"015F",X"0111",X"0103",X"0104",X"00B4",X"0074",X"0057",X"FFEF",X"FFAE",X"FF97",X"FF2A",X"FF55",X"FF45",X"FF0B",X"FF1D",X"FF2A",X"FF0B",X"FF19",X"FF07",X"FF46",X"FF9F",X"FFBF",X"FFCF",X"FF57",X"FF59",X"FF34",X"FF89",X"FF8F",X"FF7E",X"FF6D",X"FFBB",X"FFC4",X"FFC9",X"FFC4",X"FFA8",X"FFBE",X"0012",X"0037",X"005A",X"0036",X"001A",X"FFB2",X"FF4A",X"FF88",X"FF3B",X"FF4F",X"FF5D",X"FF8B",X"FFA8",X"FFB0",X"FF7F",X"FF9F",X"FF54",X"FF55",X"FF55",X"FF23",X"FF86",X"FF72",X"FF64",X"FF9A",X"FF95",X"FFD3",X"0001",X"0000",X"001C",X"003C",X"0040",X"0040",X"004D",X"FFFB",X"0066",X"0075",X"0091",X"0085",X"005C",X"FFDF",X"FFD1",X"FF9D",X"FF95",X"FFCD",X"FFA6",X"FF6C",X"FF6A",X"FF5E",X"FF9C",X"FF88",X"FF9E",X"FFEA",X"000F",X"0008",X"002A",X"0029",X"009D",X"00B7",X"010A",X"00EA",X"008A",X"0062",X"003A",X"0063",X"00E9",X"00A5",X"003D",X"0022",X"0007",X"0023",X"0088",X"0072",X"00AB",X"008D",X"FFBD",X"FFB6",X"FF93",X"0043",X"00F7",X"00E4",X"0068",X"FFE3",X"FF6F",X"FF86",X"0049",X"007A",X"00B7",X"006A",X"003A",X"FF8B",X"FFA1",X"FFDE",X"0051",X"0074",X"002E",X"FF96",X"FF94",X"FFC8",X"005E",X"00E4",X"00A8",X"004D",X"FFAA",X"FF68",X"FFDA",X"0098",X"00E0",X"00B3",X"FFEC",X"FFBC",X"001B",X"00FA",X"010D",X"00FF",X"0078",X"0039",X"003B",X"0033",X"0059",X"0073",X"0077",X"0011",X"FF9F",X"FF11",X"FF18",X"FFB6",X"0072",X"0091",X"0025",X"FF35",X"FEA2",X"FF77",X"003E",X"00F4",X"0020",X"FE91",X"FDD5",X"FEDF",X"FFE3",X"00E7",X"0002",X"FE91",X"FD97",X"FE7A",X"FFF3",X"013B",X"00E9",X"FF71",X"FDF8",X"FE09",X"FF76",X"0168",X"0210",X"00DC",X"FEDF",X"FDB6",X"FEC9",X"009A",X"01B0",X"00E0",X"FF3F",X"FD3F",X"FDCD",X"FF77",X"0155",X"0193",X"0075",X"FE47",X"FCFD",X"FDE0",X"FFD4",X"017B",X"00E3",X"FF35",X"FD14",X"FCCF",X"FECC",X"015B",X"024C",X"0128",X"FE08",X"FCB8",X"FE8E",X"0227",X"049B",X"036F",X"FFF9",X"FC8D",X"FCB2",X"007B",X"046C",X"04D2",X"0198",X"FCDF",X"FB6C",X"FEAE",X"03C4",X"0582",X"0212",X"FC38",X"F98F",X"FC0B",X"01EF",X"0574",X"0358",X"FDBF",X"F92F",X"FAC3",X"0152",X"06D8",X"0644",X"0058",X"FA6C",X"FA1D",X"FFB0",X"0689",X"07CA",X"0266",X"FAE3",X"F7D1",X"FD58",X"061D",X"09B2",X"04CE",X"FBA8",X"F656",X"FA9D",X"04F4",X"0B4B",X"0706",X"FC52",X"F440",X"F748",X"02D8",X"0BD8",X"0983",X"FDF6",X"F396",X"F434",X"FFF8",X"0B69",X"0BB8",X"00A1",X"F434",X"F255",X"FE1D",X"0B8C",X"0E91",X"034D",X"F43F",X"F082",X"FC70",X"0BFD",X"1028",X"055D",X"F5C7",X"EFCB",X"FA2A",X"0B0A",X"1292",X"0928",X"F63E",X"ED7F",X"F780",X"0A11",X"1302",X"093C",X"F578",X"EAED",X"F405",X"0771",X"1313",X"0C61",X"F81E",X"EA1D",X"F1DF",X"07E5",X"1669",X"0F6B",X"F91C",X"E891",X"EFE7",X"07A3",X"183A",X"119E",X"F8C1",X"E6F4",X"EF2B",X"08ED",X"1A57",X"1350",X"F8FB",X"E581",X"EDD9",X"0852",X"1AB3",X"12BA",X"F734",X"E4C9",X"EEBE",X"08C4",X"18A4",X"1058",X"F6E8",X"E71E",X"F184",X"09AD",X"1743",X"0DE1",X"F581",X"E716",X"F2C7",X"0B37",X"17CB",X"0BD0",X"F224",X"E5C7",X"F4D8",X"0ECC",X"193E",X"0946",X"EE66",X"E552",X"F875",X"1308",X"1A3E",X"05D0",X"E986",X"E460",X"FBCF",X"16AF",X"1A6A",X"00CC",X"E451",X"E545",X"0269",X"1C80",X"195F",X"FAE1",X"E0A2",X"E8B5",X"0A1E",X"20DD",X"1658",X"F258",X"DC8C",X"EE4A",X"1262",X"224C",X"0E16",X"E869",X"DC1E",X"F7AE",X"1BA6",X"21ED",X"0427",X"E0DB",X"E0E3",X"038C",X"2242",X"1C72",X"F7A9",X"DB71",X"E8C8",X"0FBF",X"254E",X"1238",X"EAA5",X"DB07",X"F4F6",X"1AB7",X"237B",X"04E9",X"DF45",X"DF7E",X"0482",X"2467",X"1BB3",X"F34D",X"D945",X"EC48",X"1617",X"2696",X"0A8C",X"E205",X"DD44",X"0127",X"22D5",X"1C52",X"F467",X"D9B9",X"EC6F",X"158E",X"2583",X"0956",X"E0B7",X"DD65",X"02B9",X"2413",X"1B8F",X"F171",X"D87E",X"EF48",X"1A0A",X"2758",X"0678",X"DC39",X"DEE2",X"0CC9",X"2A36",X"160B",X"E70C",X"D6E1",X"F8BD",X"2419",X"237E",X"F793",X"D557",X"E78C",X"17AE",X"2B5A",X"0957",X"DB3C",X"DAF7",X"08AA",X"2A7E",X"17CA",X"E83D",X"D74C",X"F8F3",X"2253",X"2123",X"F7AF",X"DA0B",X"ECAC",X"172D",X"244B",X"0344",X"DE48",X"E4C4",X"0D3F",X"23EB",X"0C4E",X"E3DE",X"E0F8",X"0694",X"22D6",X"11F7",X"E8EF",X"DEE9",X"007B",X"20D8",X"14C9",X"EB57",X"DC4A",X"FCCE",X"1FC4",X"17A2",X"EF56",X"DCB7",X"F87D",X"1DA3",X"1B57",X"F2A4",X"DB1F",X"F491",X"1CD6",X"1D3A",X"F3A0",X"D9A2",X"F3CB",X"1F02",X"1F5D",X"F3D9",X"D905",X"F45C",X"2035",X"1FBF",X"F358",X"D7F5",X"F4B9",X"2042",X"1F23",X"F1CE",X"D79A",X"F62C",X"20CB",X"1D0B",X"F035",X"D894",X"F8CE",X"22EF",X"1B0F",X"EC8F",X"D9A5",X"FD46",X"2467",X"1952",X"E9A5",X"DA3F",X"018F",X"2637",X"15FF",X"E63E",X"DC3D",X"0580",X"2686",X"110A",X"E2AF",X"DF09",X"0B0D",X"265A",X"09E8",X"DF55",X"E5CA",X"1233",X"23BA",X"009D",X"DDA4",X"EEB1",X"18E5",X"1D0F",X"F617",X"DF57",X"FA40",X"1D73",X"14CE",X"EB70",X"E253",X"05F4",X"2160",X"0989",X"E202",X"E861",X"11BF",X"2083",X"FDC2",X"DDFA",X"F222",X"1ABA",X"1A2A",X"F10D",X"E0BE",X"00C3",X"1F5A",X"0BF1",X"E6ED",X"EAFF",X"0FBA",X"1AC1",X"F98F",X"E48A",X"FC3D",X"19D0",X"0D28",X"E9E2",X"E99D",X"0D3B",X"1AE9",X"FBB4",X"E461",X"FA80",X"18DC",X"0E5E",X"EE04",X"EF06",X"0D08",X"14A9",X"F8F5",X"ECD3",X"03E6",X"1441",X"0136",X"EC03",X"FAF6",X"1395",X"0ABA",X"EEF9",X"F167",X"0E0A",X"1323",X"F578",X"EAD0",X"066F",X"1885",X"FF2C",X"E5F4",X"FA7E",X"1B6C",X"0EA0",X"E5F0",X"E94F",X"13F3",X"1E99",X"F561",X"DD8B",X"FFBD",X"2213",X"0A4C",X"DF88",X"EC90",X"1884",X"1949",X"ED57",X"E154",X"092C",X"1EB3",X"FDDE",X"E13B",X"F963",X"1C6D",X"0C91",X"E682",X"EE03",X"144F",X"1655",X"F05D",X"E75C",X"07DF",X"1988",X"FBD0",X"E539",X"FC8C",X"1809",X"0616",X"E78E",X"F55B",X"14E3",X"0DB5",X"EBDA",X"EED9",X"1157",X"157C",X"F184",X"E6D6",X"09F7",X"1D95",X"FC39",X"E0C0",X"FD42",X"1E79",X"09E2",X"E414",X"F11E",X"178F",X"14BE",X"EB2A",X"E7E0",X"1063",X"1C6F",X"F576",X"E2CB",X"04F7",X"1EF5",X"01D0",X"E043",X"F83D",X"1E14",X"0E19",X"E4AF",X"EE7C",X"17D5",X"181B",X"EBB7",X"E4CA",X"0ED1",X"1E06",X"F424",X"DEC2",X"0472",X"21D1",X"0063",X"DCBE",X"F874",X"216A",X"0E11",X"E11D",X"EE79",X"1C10",X"17B2",X"E7F8",X"E646",X"1461",X"1E3F",X"EFA3",X"E04B",X"0AC9",X"2221",X"FA95",X"DC65",X"FEAB",X"22BA",X"05E0",X"DDD6",X"F4D4",X"1EDC",X"0F07",X"E2CF",X"EE22",X"19B4",X"154C",X"E815",X"E88E",X"14FF",X"1B75",X"ED61",X"E273",X"0CEE",X"20A3",X"F74A",X"DF33",X"044E",X"2302",X"01BB",X"E01B",X"FC04",X"20F1",X"0B0D",X"E171",X"F1DE",X"1CE5",X"13F5",X"E60B",X"EA13",X"1677",X"18DF",X"EBE2",X"E650",X"100C",X"1C00",X"F20B",X"E22C",X"08B6",X"1EEB",X"F89D",X"DF15",X"0191",X"2119",X"0149",X"DE37",X"FAE3",X"213E",X"08B4",X"E023",X"F4A6",X"1ED2",X"102F",X"E3E3",X"EDA5",X"1A4F",X"1741",X"E7F6",X"E7B5",X"1449",X"19EA",X"EDE9",X"E5C6",X"0DE5",X"1B2C",X"F2D6",X"E3C1",X"088D",X"1D43",X"F847",X"E05A",X"03B1",X"2039",X"FEA2",X"DE1B",X"FCB1",X"1FAE",X"05DF",X"E0BB",X"F722",X"1C63",X"0B9C",X"E565",X"F2AD",X"1950",X"10EB",X"E838",X"EE50",X"1584",X"1312",X"EC0C",X"ECB6",X"1203",X"137F",X"ED45",X"EB51",X"1038",X"1599",X"EF99",X"E760",X"0C03",X"1947",X"F44A",X"E3E0",X"07FC",X"1B21",X"F8A7",X"E511",X"0571",X"1A9E",X"FB94",X"E3A6",X"0186",X"1CFB",X"0031",X"E236",X"FD62",X"1E53",X"0756",X"E3EA",X"F8C1",X"1D27",X"0BC6",X"E4A7",X"F429",X"1B1E",X"1015",X"E590",X"EDFE",X"1840",X"152F",X"E821",X"E8C9",X"1441",X"1A1D",X"EE06",X"E63F",X"1006",X"1BAF",X"F1A2",X"E341",X"0A66",X"1DBB",X"F698",X"E02C",X"04D6",X"2093",X"FCBC",X"DF0C",X"FF85",X"2059",X"03AD",X"DF89",X"F92A",X"1FD5",X"09FD",X"E043",X"F442",X"203E",X"0F18",X"E14F",X"EF57",X"1D46",X"135C",X"E426",X"EBC2",X"1963",X"1664",X"E859",X"E8C3",X"155B",X"18D1",X"EC22",X"E6EF",X"126D",X"1B3E",X"EF7C",X"E559",X"0FE7",X"1CD2",X"F441",X"E3FC",X"0A12",X"1E09",X"F91C",X"E2CB",X"0526",X"1DF8",X"FD7B",X"E431",X"03A7",X"1DC4",X"FF80",X"E44E",X"00EF",X"1D34",X"016E",X"E2D0",X"FCD4",X"1C0A",X"03A4",X"E27D",X"F909",X"1B54",X"07E4",X"E3B6",X"F58A",X"1AE8",X"0B09",X"E455",X"F236",X"1957",X"0E3E",X"E52C",X"EFD0",X"1870",X"1088",X"E64C",X"ED8E",X"16D8",X"11C7",X"E85F",X"EBF2",X"1490",X"14BC",X"EAE4",X"E930",X"11AA",X"1767",X"EE03",X"E6C9",X"0FD7",X"1A0D",X"F217",X"E644",X"0C42",X"1A1A",X"F485",X"E53C",X"093F",X"1B98",X"F75B",X"E460",X"0648",X"1D8A",X"FC93",X"E340",X"0249",X"1D96",X"0015",X"E2FC",X"FEE3",X"1E88",X"036E",X"E191",X"FC4A",X"1F73",X"0776",X"E36F",X"F726",X"1C2A",X"0C45",X"E4A6",X"F0D4",X"17E4",X"0FBC",X"E6B8",X"EBB3",X"142B",X"133D",X"E82E",X"E787",X"11C9",X"16BA",X"EB8B",X"E3DA",X"0DD5",X"1B28",X"F2BC",X"E4B5",X"0AFD",X"1DE7",X"F9A8",X"E53E",X"06FC",X"1EC1",X"FE4B",X"E41A",X"02BE",X"1DFA",X"0170",X"E3B9",X"FE31",X"1D3A",X"05DF",X"E460",X"F9B4",X"1BD3",X"0A2A",X"E591",X"F3EF",X"1A39",X"0EC8",X"E602",X"EE64",X"183F",X"1408",X"E7E5",X"EAAF",X"1622",X"17D2",X"EC2A",X"E79B",X"1135",X"1953",X"F01C",X"E648",X"0D9E",X"1AD9",X"F4EA",X"E566",X"09A3",X"1C38",X"F92E",X"E46F",X"04BC",X"1CD0",X"FDC6",X"E38F",X"FFAC",X"1D0A",X"02BF",X"E392",X"FAE7",X"1BD0",X"0834",X"E4EE",X"F596",X"197E",X"0D02",X"E6E9",X"F0F9",X"15E3",X"0FDE",X"EB33",X"EE52",X"129C",X"13C9",X"EDE2",X"EC56",X"105E",X"1552",X"F240",X"EA72",X"0C69",X"18E4",X"F672",X"E7ED",X"07DA",X"18BF",X"F9D9",X"E6B4",X"0429",X"1983",X"FE83",X"E6A6",X"FFF0",X"1A8B",X"0379",X"E6B7",X"FB02",X"1A08",X"07B9",X"E782",X"F788",X"18DD",X"0BC2",X"E7F8",X"F319",X"172E",X"0FF2",X"E9B3",X"EF13",X"142D",X"114F",X"EABC",X"EB7D",X"0FE2",X"13C4",X"EDC7",X"E820",X"0C45",X"176E",X"F1D5",X"E552",X"08E4",X"19B3",X"F7FE",X"E54F",X"0536",X"1B55",X"FDC3",X"E575",X"00BE",X"1B7E",X"02E2",X"E3FF",X"F942",X"186C",X"0664",X"E4BA",X"F4F2",X"1749",X"0C13",X"E7C9",X"F0D2",X"1482",X"10F7",X"EC13",X"EDE8",X"11B5",X"15C1",X"F222",X"EB9A",X"0E70",X"19DF",X"F5F5",X"E6D1",X"078B",X"18A8",X"F7FD",X"E4A1",X"0310",X"19F5",X"001D",X"E77D",X"FF8F",X"19E7",X"02F6",X"E5E4",X"F994",X"1845",X"075C",X"E6B0",X"F6E3",X"19C6",X"0E0A",X"EA2F",X"F351",X"164F",X"10DB",X"ED42",X"EE41",X"0F7B",X"11FE",X"F17F",X"ED59",X"0E17",X"16A2",X"F579",X"EAC4",X"0AC8",X"1788",X"F647",X"E76D",X"07A4",X"19D1",X"FC7C",X"E97D",X"067F",X"1D34",X"0197",X"E974",X"0177",X"19D9",X"0294",X"E6D7",X"F87E",X"156D",X"0774",X"E75C",X"F397",X"1559",X"0D91",X"E97A",X"EF03",X"0FCE",X"0E8E",X"EC6B",X"EAEC",X"0E0E",X"14DF",X"F302",X"EBD3",X"0CFB",X"1945",X"F77F",X"E7E8",X"0631",X"1794",X"FA3D",X"E4A3",X"0039",X"1911",X"0057",X"E5DB",X"FE21",X"1A10",X"0322",X"E4A0",X"F7E0",X"1652",X"068E",X"E606",X"F47F",X"15A1",X"0E15",X"EBB1",X"F063",X"12E8",X"12BF",X"EE19",X"EB7A",X"0E24",X"13B2",X"F03A",X"E910",X"0A8B",X"17AC",X"F7EE",X"E856",X"061D",X"18C9",X"FA5E",X"E39E",X"FF76",X"17D3",X"010A",X"E8C8",X"FCDF",X"19EC",X"099D",X"E8FC",X"F773",X"1825",X"0B7E",X"E7BC",X"F27D",X"1561",X"0E77",X"EB19",X"EFC5",X"124C",X"1300",X"EEA9",X"EB33",X"0D3C",X"156D",X"F2E9",X"E8DB",X"0A6A",X"1A15",X"FABD",X"E936",X"07D4",X"1B58",X"FEDE",X"E7EE",X"00DB",X"19BF",X"021E",X"E634",X"FAE9",X"17F2",X"0732",X"E942",X"F8DE",X"1766",X"0BDF",X"EA55",X"F2DC",X"13AC",X"0E72",X"ED7A",X"EFDC",X"1238",X"148B",X"F266",X"ED24",X"0D5E",X"15DD",X"F3AF",X"E7D7",X"065D",X"143A",X"F711",X"E703",X"0267",X"16A6",X"FE84",X"E7D4",X"FF2E",X"1800",X"0272",X"E7FA",X"FACC",X"1692",X"0681",X"EA33",X"FA28",X"1763",X"0DEB",X"EE52",X"F51E",X"1563",X"10E9",X"ED88",X"EFD5",X"1114",X"1144",X"EFE4",X"EDB3",X"0D4B",X"13BE",X"F454",X"EBD8",X"0A5A",X"14DA",X"F7D7",X"EA62",X"0633",X"166B",X"FEB9",X"EC03",X"03A2",X"18BD",X"0228",X"EAA1",X"FE9A",X"152F",X"03E8",X"E950",X"F7E4",X"11F1",X"06CF",X"EC13",X"F721",X"124D",X"0BCA",X"EF1D",X"F2C0",X"0FE2",X"0DB7",X"F0CC",X"F06F",X"0D56",X"116E",X"F2DF",X"EDB5",X"0A9B",X"12D6",X"F63B",X"EB71",X"0738",X"1350",X"F792",X"E948",X"03B2",X"131A",X"FC92",X"EBA8",X"012F",X"1546",X"00F5",X"EA9A",X"FDB0",X"1419",X"03E4",X"EC8E",X"FC64",X"136C",X"0726",X"EE65",X"F8A9",X"1259",X"09C0",X"EF1D",X"F738",X"0F91",X"092F",X"EE53",X"F1F5",X"0B5C",X"0AE6",X"F1DD",X"F1BC",X"0BE9",X"0E16",X"F63A",X"F159",X"0A52",X"111B",X"F99D",X"F0C9",X"059C",X"108A",X"FBCA",X"EE6C",X"03FF",X"11B7",X"FD11",X"EE12",X"00D8",X"102B",X"FC0E",X"EC0C",X"FE59",X"11D5",X"0254",X"EF50",X"FDB5",X"1257",X"05F6",X"EFDD",X"FBD7",X"1075",X"06AB",X"F059",X"F7E3",X"0E8C",X"083D",X"F1E8",X"F7A9",X"0D71",X"0AC4",X"F32C",X"F354",X"09B4",X"0B21",X"F3C8",X"F1FA",X"0948",X"0D2A",X"F73B",X"F216",X"08DB",X"1011",X"FB40",X"F1AA",X"058B",X"0FEC",X"FB5E",X"EFBB",X"0397",X"0FD2",X"FEA3",X"F1BD",X"01EF",X"0F29",X"FF5A",X"F010",X"FDC6",X"0C5E",X"00B1",X"F1AA",X"FC3D",X"0C39",X"0381",X"F202",X"FC51",X"0D8E",X"05CA",X"F3D0",X"FB1F",X"0BFB",X"053A",X"F416",X"F8EC",X"09C8",X"073E",X"F554",X"F80F",X"09A6",X"079D",X"F747",X"F8D0",X"095E",X"094D",X"F8FB",X"F7FF",X"07D8",X"09CC",X"FA75",X"F712",X"0691",X"0B33",X"FB0D",X"F649",X"0574",X"0B96",X"FCF6",X"F528",X"02CD",X"0B7A",X"FE27",X"F4FB",X"01D4",X"0BED",X"0037",X"F617",X"014C",X"0CE5",X"00B6",X"F3EA",X"FDDB",X"0BAA",X"02AC",X"F4A7",X"FE9A",X"0C74",X"04F3",X"F5AC",X"FC1B",X"0A5A",X"040D",X"F406",X"F829",X"07E9",X"051A",X"F596",X"F847",X"06EE",X"0834",X"F774",X"F640",X"060F",X"066A",X"F760",X"F4F6",X"0586",X"0A6B",X"FBE7",X"F79C",X"06C9",X"0C1D",X"FC09",X"F475",X"0247",X"08EB",X"FB55",X"F287",X"0128",X"0CD8",X"0178",X"F420",X"006D",X"0E4B",X"02D7",X"F387",X"FB4D",X"0A67",X"03B4",X"F413",X"FAAE",X"0AB2",X"06BE",X"F631",X"F90A",X"0865",X"069A",X"F4A9",X"F405",X"0536",X"06E0",X"F741",X"F523",X"060F",X"0A69",X"FAD8",X"F4B3",X"033D",X"0B11",X"FBEB",X"F264",X"01A6",X"0BE5",X"FED1",X"F4CC",X"029D",X"0C52",X"0026",X"F506",X"FFF0",X"0C71",X"0183",X"F33D",X"FCEB",X"0C05",X"0598",X"F4FF",X"FC8F",X"0BEB",X"0573",X"F4B4",X"F922",X"095D",X"05CF",X"F5F6",X"FAC0",X"0B4B",X"090D",X"F825",X"F9BC",X"0A4A",X"0A1E",X"F95A",X"F73A",X"0757",X"091B",X"FA30",X"F6D0",X"0889",X"0CBD",X"FD76",X"F81A",X"06BD",X"0D00",X"FCEB",X"F3E3",X"0367",X"0C94",X"FF02",X"F46C",X"00A5",X"0C03",X"FFE6",X"F36A",X"FE5C",X"09C9",X"FFC2",X"F363",X"FC65",X"0ADB",X"02F9",X"F5B3",X"FD77",X"0C26",X"055F",X"F63D",X"FB32",X"09B1",X"051F",X"F62D",X"F8A0",X"092D",X"07D7",X"F630",X"F743",X"08CB",X"08FB",X"F876",X"F63D",X"067C",X"092D",X"F996",X"F4F0",X"044D",X"0AAB",X"FD14",X"F58E",X"02DD",X"0A02",X"FBF6",X"F37F",X"FFD2",X"08D6",X"FE78",X"F49D",X"FFE2",X"09CF",X"0003",X"F593",X"FEA2",X"0A03",X"0348",X"F724",X"FC83",X"079A",X"02BA",X"F6E9",X"FBC5",X"094A",X"07E0",X"F8ED",X"F96D",X"0732",X"069C",X"F8CB",X"F776",X"05A4",X"08B2",X"FB54",X"F6A0",X"013C",X"062E",X"FBA7",X"F4E2",X"003E",X"07E9",X"FDFA",X"F4C8",X"FD72",X"067F",X"007A",X"F6B6",X"FE76",X"09B1",X"027F",X"F756",X"FC68",X"0796",X"0370",X"F6F2",X"FAD4",X"0892",X"05B8",X"F6EF",X"F881",X"077C",X"07EF",X"F9D4",X"F98B",X"07C4",X"079B",X"F96D",X"F7ED",X"061F",X"09B8",X"FD5F",X"F9D1",X"0473",X"08B2",X"FC1A",X"F62A",X"0342",X"0825",X"FC57",X"F7AB",X"0382",X"092D",X"FD06",X"F572",X"01B2",X"0C58",X"0175",X"F749",X"0103",X"0A8F",X"0222",X"F717",X"003B",X"0C62",X"0557",X"F8BA",X"FC89",X"09C8",X"0602",X"F926",X"FE0A",X"09EA",X"066A",X"F925",X"FAAD",X"06B2",X"0454",X"F881",X"FA08",X"06B3",X"072F",X"FA28",X"F6E0",X"0344",X"06D5",X"FA89",X"F7B5",X"052B",X"0B12",X"FCA5",X"F593",X"01F0",X"090C",X"0077",X"F854",X"00DD",X"09BF",X"0135",X"F702",X"FE17",X"07C7",X"014A",X"F7BB",X"FF98",X"09EB",X"02D1",X"F50D",X"FAF9",X"07AE",X"0353",X"F64A",X"F9F1",X"0751",X"0411",X"F574",X"F7B0",X"07A7",X"0801",X"F80B",X"F578",X"0287",X"04C2",X"F7F1",X"F4FD",X"0357",X"083F",X"FC37",X"F79F",X"03F8",X"08D3",X"FBF3",X"F591",X"011E",X"097D",X"FE6F",X"F688",X"00E3",X"098A",X"FE74",X"F56D",X"0002",X"0B96",X"033B",X"F597",X"FBB0",X"0827",X"0294",X"F677",X"FBCA",X"0947",X"052A",X"F5F1",X"FA04",X"07D4",X"0513",X"F65F",X"F847",X"06D5",X"0548",X"F7F1",X"F900",X"06EC",X"071F",X"F95A",X"F7C1",X"0674",X"08D8",X"FB18",X"F570",X"0297",X"08BC",X"FDA5",X"F804",X"048E",X"0AAC",X"FE54",X"F626",X"0265",X"0C95",X"017F",X"F63F",X"FF7C",X"0982",X"00FE",X"F5CE",X"FF15",X"0ABC",X"0293",X"F6FF",X"FD40",X"0889",X"035F",X"F739",X"FAE2",X"06F5",X"042D",X"FA62",X"FD07",X"06DD",X"0398",X"F707",X"FA8B",X"0804",X"07EB",X"FB95",X"F9A1",X"0537",X"0894",X"FCA6",X"FA7B",X"05B1",X"08D4",X"FDA6",X"F84E",X"030E",X"08B2",X"FF76",X"F950",X"00E3",X"075B",X"FF9A",X"FA0B",X"040C",X"086B",X"FE26",X"F81A",X"00D8",X"07C1",X"FF72",X"F67E",X"FE9D",X"072C",X"0195",X"F8F1",X"FE37",X"07A8",X"037C",X"FA11",X"FD46",X"061C",X"038B",X"FA4B",X"FB70",X"0552",X"044D",X"FA3D",X"FAAB",X"054A",X"06ED",X"FC32",X"F8F5",X"032B",X"0543",X"FBA9",X"F8D0",X"0262",X"063C",X"FCFC",X"F7B3",X"FF82",X"0534",X"FEBE",X"F96A",X"01AE",X"07DF",X"00B0",X"F9AE",X"00C2",X"0875",X"022C",X"F8B5",X"FDF2",X"0814",X"0430",X"F963",X"FAD5",X"0410",X"0175",X"F89F",X"FBB1",X"0567",X"0465",X"FA52",X"FB07",X"0445",X"0396",X"FA12",X"F9F9",X"03A1",X"04F8",X"FC08",X"F99A",X"0362",X"065C",X"FDA8",X"F9EE",X"02F6",X"073B",X"FE8A",X"F90E",X"003F",X"0411",X"FC03",X"F6EE",X"001A",X"0660",X"FE37",X"F638",X"FDDA",X"079A",X"026F",X"F923",X"FE87",X"074D",X"024B",X"F91C",X"FDC1",X"0718",X"0222",X"F86C",X"FC63",X"072B",X"04EB",X"F9BF",X"FB55",X"0667",X"0575",X"F8AB",X"F7E5",X"03AF",X"0630",X"FC35",X"F90A",X"01E8",X"0539",X"FC7C",X"F816",X"0142",X"07E7",X"002F",X"FA53",X"014C",X"0674",X"FF0A",X"F896",X"FFD6",X"074D",X"0168",X"FA59",X"0006",X"0894",X"03E0",X"F9C0",X"FC31",X"072F",X"076A",X"FF56",X"FF44",X"06EF",X"05A2",X"FD07",X"FD32",X"056A",X"04D3",X"FD50",X"FD66",X"068E",X"0743",X"FDE5",X"FA1F",X"02B5",X"068A",X"FF5F",X"FAFF",X"028B",X"0706",X"FF0A",X"F9F0",X"0097",X"05B7",X"FFC6",X"FB32",X"01F5",X"06D0",X"FF27",X"F90A",X"FF67",X"0629",X"FFBA",X"F826",X"FCF5",X"0375",X"FE8B",X"F98B",X"FFDB",X"063D",X"FF82",X"F81F",X"FD02",X"0427",X"005F",X"F9D4",X"FEB8",X"06CE",X"0333",X"FB2F",X"FEA9",X"0592",X"01F9",X"F999",X"FC89",X"0593",X"030D",X"FA17",X"FC08",X"04D4",X"02AB",X"F9AD",X"FA48",X"0278",X"027F",X"FB08",X"FBDB",X"0503",X"047B",X"FA76",X"F95F",X"0267",X"03A0",X"FB86",X"FACD",X"044E",X"0622",X"FDA2",X"F9D1",X"0058",X"02BB",X"FBDA",X"FAE1",X"02C2",X"056F",X"FE06",X"FA28",X"0083",X"03D0",X"FD28",X"F9A7",X"FFF2",X"04CB",X"00BF",X"FD4C",X"01A6",X"044E",X"FEB3",X"FA7E",X"FF70",X"05CC",X"0200",X"FBFE",X"FFA7",X"0453",X"0090",X"FBB3",X"FFA2",X"0559",X"02C9",X"FC0B",X"FDE8",X"045B",X"034F",X"FE09",X"FF2C",X"0330",X"00DC",X"FC01",X"FD6D",X"0362",X"0354",X"FD3E",X"FCAE",X"038E",X"04F2",X"FF2B",X"FCDE",X"010B",X"02C6",X"FDAE",X"FBB7",X"00F5",X"03E9",X"FF40",X"FBD0",X"FF83",X"01A9",X"FD53",X"FBED",X"015F",X"0434",X"FF04",X"FB45",X"FF4A",X"037F",X"FF63",X"FB1A",X"FEAC",X"0367",X"0043",X"FB82",X"FE9A",X"03EE",X"021E",X"FD01",X"FEB6",X"0404",X"01D6",X"FC84",X"FED6",X"0471",X"0381",X"FF71",X"00AF",X"0501",X"03C4",X"FEB3",X"FEA9",X"03AB",X"0477",X"FEE0",X"FCF1",X"01B9",X"0379",X"FF87",X"FE0C",X"0261",X"041A",X"FEF1",X"FC7C",X"00E3",X"03A8",X"FF7D",X"FCEA",X"00CC",X"03BD",X"00A1",X"FE0E",X"002F",X"0267",X"FFC4",X"FC49",X"FE9C",X"029F",X"00D9",X"FD02",X"FEDA",X"02BF",X"0051",X"FC47",X"FDB3",X"01BA",X"013E",X"FD49",X"FD73",X"0192",X"01F8",X"FE21",X"FD5B",X"00A9",X"0129",X"FD72",X"FC61",X"FFB4",X"0145",X"FEAC",X"FDF0",X"00EA",X"02AC",X"FFF0",X"FEB0",X"01FF",X"03C4",X"FFDA",X"FD54",X"006F",X"032B",X"003F",X"FD4F",X"FEB8",X"00A4",X"FF4F",X"FD36",X"FEDF",X"0160",X"FF90",X"FC22",X"FC74",X"FF5E",X"002D",X"FE51",X"FF28",X"023B",X"01E7",X"FEC0",X"FF58",X"02C9",X"032A",X"FFAC",X"FE71",X"FF70",X"FF4A",X"FDDD",X"FDF8",X"FFEF",X"FFE3",X"FD29",X"FC1B",X"FF06",X"00EF",X"FF4C",X"FE46",X"00AC",X"01E3",X"FFB1",X"FE0B",X"FEDF",X"0026",X"FF3A",X"FDE4",X"FF32",X"00BB",X"FFB2",X"FD62",X"FD78",X"FFA7",X"005F",X"FFF5",X"00FC",X"0256",X"01F2",X"00F5",X"013F",X"022D",X"0125",X"FF69",X"010E",X"024B",X"022B",X"0137",X"00F4",X"014E",X"0120",X"FFC9",X"FEFF",X"007A",X"01C5",X"00B3",X"FF35",X"FF48",X"FF75",X"FEB3",X"FE5A",X"FFB4",X"00D6",X"0090",X"0063",X"0166",X"025B",X"01BE",X"FFE1",X"FF18",X"FF61",X"FEE0",X"FE5B",X"FF6A",X"00BB",X"006D",X"FF42",X"FF57",X"009C",X"0106",X"FFEF",X"FFC3",X"0088",X"00F1",X"0028",X"0004",X"008E",X"0040",X"FF65",X"FF34",X"003F",X"0111",X"006A",X"FFE8",X"000B",X"0014",X"FF30",X"FF09",X"FFF3",X"0079",X"0017",X"FF72",X"FF56",X"0017",X"005A",X"00AE",X"00EE",X"00BF",X"FFF9",X"FFAC",X"0077",X"010A",X"0083",X"FFAF",X"FFDB",X"0040",X"0043",X"FF77",X"FF81",X"FFDF",X"FFFF",X"FFEC",X"0072",X"0124",X"0103",X"0091",X"0096",X"0134",X"0191",X"00F8",X"00A8",X"00ED",X"00E8",X"0061",X"FFF3",X"FFC4",X"FF26",X"FEDF",X"FF08",X"FF94",X"0031",X"007E",X"00E9",X"00C5",X"0040",X"FF7A",X"FED4",X"FEC5",X"FFD2",X"0132",X"0107",X"FFD7",X"FF5B",X"FF8E",X"FF75",X"FF19",X"FF0B",X"FF51",X"003A",X"007A",X"FFF5",X"FF23",X"FF1B",X"FF11",X"FF2E",X"FF8A",X"FF53",X"FF2D",X"FF6B",X"FF48",X"FF1E",X"FEE7",X"FEA9",X"FE88",X"FECB",X"FF43",X"FEE4",X"FE53",X"FE9D",X"FF1A",X"FF59",X"FF0C",X"FEA4",X"FE88",X"FEF4",X"FF61",X"FF81",X"FF88",X"FFD1",X"FFDB",X"00B3",X"01BC",X"0231",X"0180",X"0096",X"0003",X"FF7B",X"FF03",X"FF13",X"FFF1",X"FFFE",X"FFB6",X"FF67",X"FF39",X"FF2B",X"FF4D",X"FFE0",X"0072",X"0060",X"FF8C",X"FF00",X"FFA7",X"007A",X"00DC",X"0088",X"0042",X"0053",X"0069",X"009E",X"0096",X"0066",X"000E",X"FFE5",X"0001",X"005C",X"0007",X"FFA5",X"001F",X"00E1",X"00CD",X"006F",X"00B8",X"017C",X"019D",X"00FC",X"008D",X"0079",X"004B",X"005F",X"00C4",X"0100",X"0045",X"FF24",X"FF1C",X"FFED",X"FFF0",X"FEE6",X"FEAA",X"FF25",X"FFB6",X"0001",X"FFFA",X"0065",X"0094",X"0066",X"001E",X"006A",X"011E",X"0167",X"00D2",X"010A",X"0160",X"0103",X"0038",X"FFDD",X"002C",X"FFEE",X"FF38",X"FEE3",X"FEC0",X"FE5F",X"FE1F",X"FE84",X"FF12",X"FF5B",X"FF46",X"FFB5",X"0083",X"009D",X"005E",X"0066",X"00D3",X"00F3",X"0097",X"0004",X"FF54",X"FF96",X"FF84",X"FF55",X"FFDB",X"0074",X"002C",X"FF72",X"FF76",X"0020",X"0099",X"0076",X"0072",X"00A4",X"00C3",X"0101",X"0096",X"00BF",X"0119",X"00CF",X"00B4",X"00C5",X"00E8",X"0065",X"FFCE",X"FF68",X"FF2B",X"FF3B",X"FF36",X"FF80",X"FF9E",X"FF45",X"FECC",X"FF50",X"0043",X"0081",X"0047",X"009B",X"01D0",X"01CC",X"00E0",X"004F",X"0053",X"0031",X"FF7F",X"FEDF",X"FE36",X"FDE3",X"FE3E",X"FEC3",X"FF67",X"FF86",X"FF7D",X"FF9B",X"0000",X"FFF4",X"FF52",X"FEDB",X"FF31",X"FFC2",X"0087",X"0118",X"00FD",X"009E",X"002D",X"FFE5",X"FFBD",X"FFA0",X"FEBC",X"FDC3",X"FE04",X"FEDD",X"FF8F",X"FFF9",X"00BB",X"014A",X"0131",X"010F",X"00D3",X"010E",X"00C0",X"004A",X"FFFC",X"001F",X"0051",X"006B",X"0082",X"00E4",X"00EF",X"00A3",X"0074",X"0062",X"0014",X"FFCE",X"FF9B",X"FFB1",X"FFD5",X"FF77",X"FF95",X"001E",X"00E0",X"00DC",X"0087",X"00BD",X"0136",X"0125",X"0079",X"FFF0",X"FF1F",X"FEA4",X"FE70",X"FEC6",X"FF31",X"FFC0",X"0068",X"00EE",X"00DC",X"007E");
begin
 
   
 process(resetN, CLK)
	 type noteArrd is array (0 to 12) of integer;
	 variable dataTmp : noteArrd;
 begin
	if (resetN='0') then
		dataTmp := (others  => 0);
	elsif(rising_edge(CLK)) then
		dataTmp := (others  => 0);
		for i in 0 to 12 loop
			if addrArr(i) < array_size then
				if conv_integer(addrArr(i)) > 0 then
					dataTmp(i) := conv_integer(sound0(conv_integer(addrArr(i))));
				end if;
			else
				dataTmp(i) := 0;
			end if;
		end loop;
	end if;
	Q <= conv_std_logic_vector(dataTmp(0) + dataTmp(1) + dataTmp(2) + dataTmp(3) + dataTmp(4) + dataTmp(5) + dataTmp(6) + dataTmp(7) + dataTmp(8) + dataTmp(9) + dataTmp(10) + dataTmp(11) + dataTmp(12), 16);
end process;
	 

		   
end arch;